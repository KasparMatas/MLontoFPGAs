`timescale 1ns / 1ps

`define CLOCK 20 
`define DATA_WIDTH 16
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02.03.2019 16:05:53
// Design Name: 
// Module Name: first_cell_check
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module generated_model_simulator();

event error;
always @ (error) begin
    $display("ERROR at time %t", $time);
    #`CLOCK $stop;
end

task check_output(input [`DATA_WIDTH*4-1:0] result, input [`DATA_WIDTH*4-1:0] golden);
begin
    if (result!=golden) begin
        $display("Output is %0d which should be %0d instead!", result, golden);
        //->error;
    end
end
endtask

reg[31:0] file_lines_read;
integer data_file;
reg[31:0] captured_data;
reg[7:0] pixel_data [0:1023];
reg[9:0] pixels_fed;
reg[7:0] numbers_streamed;

task open_data_file(input [1023:0] file_name);
begin
  data_file = $fopen(file_name, "r");
  if (data_file == 0) begin
    $display("File %s handle was NULL", file_name);
    $stop;
  end
  else begin 
    file_lines_read = 0;
    while (!$feof(data_file)) begin
      $fscanf(data_file, "%d\n", captured_data); 
      pixel_data[file_lines_read] = captured_data;
      file_lines_read = file_lines_read + 1;
    end
  end
end
endtask

reg clk;

wire [`DATA_WIDTH*4:0] ground;
assign ground = 0;
reg [10-1:0] input_index;
reg [`DATA_WIDTH-1:0] input_value;
reg input_enable;
wire [10-1:0] index_0_0_1;
wire [`DATA_WIDTH-1:0] value_0_0_1;
wire [`DATA_WIDTH*4:0] result_0_0_1;
wire enable_0_0_1;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd91, 8'd82, 8'd145, 8'd103, 8'd69, 8'd128, 8'd62, 8'd144, 8'd42, 8'd111, 8'd45, 8'd84, 8'd114, 8'd118, 8'd96, 8'd145, 8'd150, 8'd72, 8'd109, 8'd102, 8'd61, 8'd79, 8'd144, 8'd130, 8'd148, 8'd80, 8'd135, 8'd164, 8'd167, 8'd159, 8'd113, 8'd74, 8'd115, 8'd105, 8'd70, 8'd119, 8'd110, 8'd87, 8'd125, 8'd46, 8'd103, 8'd67, 8'd119, 8'd77, 8'd50, 8'd82, 8'd89, 8'd127, 8'd109, 8'd149, 8'd152, 8'd169, 8'd150, 8'd113, 8'd109, 8'd80, 8'd77, 8'd80, 8'd71, 8'd134, 8'd133, 8'd88, 8'd84, 8'd99, 8'd92, 8'd69, 8'd149, 8'd121, 8'd93, 8'd74, 8'd97, 8'd110, 8'd80, 8'd78, 8'd139, 8'd110, 8'd101, 8'd106, 8'd111, 8'd105, 8'd152, 8'd95, 8'd110, 8'd79, 8'd93, 8'd141, 8'd156, 8'd145, 8'd146, 8'd96, 8'd80, 8'd116, 8'd167, 8'd146, 8'd145, 8'd109, 8'd150, 8'd155, 8'd105, 8'd90, 8'd136, 8'd170, 8'd111, 8'd147, 8'd87, 8'd142, 8'd86, 8'd124, 8'd142, 8'd169, 8'd132, 8'd84, 8'd133, 8'd96, 8'd153, 8'd114, 8'd149, 8'd90, 8'd109, 8'd164, 8'd129, 8'd141, 8'd101, 8'd69, 8'd112, 8'd105, 8'd99, 8'd90, 8'd148, 8'd98, 8'd157, 8'd81, 8'd141, 8'd62, 8'd109, 8'd142, 8'd141, 8'd155, 8'd146, 8'd114, 8'd126, 8'd118, 8'd83, 8'd139, 8'd147, 8'd169, 8'd127, 8'd155, 8'd127, 8'd154, 8'd167, 8'd120, 8'd150, 8'd150, 8'd79, 8'd151, 8'd112, 8'd148, 8'd79, 8'd78, 8'd139, 8'd97, 8'd105, 8'd150, 8'd130, 8'd128, 8'd117, 8'd166, 8'd89, 8'd74, 8'd122, 8'd106, 8'd128, 8'd140, 8'd95, 8'd137, 8'd126, 8'd185, 8'd140, 8'd130, 8'd153, 8'd168, 8'd167, 8'd149, 8'd127, 8'd112, 8'd116, 8'd148, 8'd159, 8'd100, 8'd127, 8'd143, 8'd149, 8'd112, 8'd130, 8'd127, 8'd83, 8'd97, 8'd129, 8'd82, 8'd117, 8'd173, 8'd102, 8'd162, 8'd180, 8'd135, 8'd164, 8'd177, 8'd128, 8'd147, 8'd66, 8'd151, 8'd72, 8'd67, 8'd170, 8'd105, 8'd99, 8'd95, 8'd135, 8'd137, 8'd191, 8'd151, 8'd126, 8'd164, 8'd130, 8'd103, 8'd94, 8'd128, 8'd161, 8'd128, 8'd154, 8'd100, 8'd107, 8'd128, 8'd116, 8'd170, 8'd175, 8'd145, 8'd151, 8'd121, 8'd122, 8'd69, 8'd89, 8'd108, 8'd97, 8'd127, 8'd120, 8'd126, 8'd200, 8'd83, 8'd156, 8'd104, 8'd102, 8'd137, 8'd91, 8'd171, 8'd170, 8'd179, 8'd158, 8'd133, 8'd180, 8'd185, 8'd166, 8'd168, 8'd134, 8'd71, 8'd97, 8'd150, 8'd118, 8'd163, 8'd75, 8'd79, 8'd162, 8'd156, 8'd83, 8'd118, 8'd153, 8'd155, 8'd115, 8'd74, 8'd70, 8'd139, 8'd83, 8'd99, 8'd99, 8'd97, 8'd172, 8'd151, 8'd99, 8'd149, 8'd180, 8'd165, 8'd117, 8'd91, 8'd66, 8'd125, 8'd136, 8'd115, 8'd159, 8'd147, 8'd86, 8'd120, 8'd145, 8'd113, 8'd122, 8'd92, 8'd86, 8'd76, 8'd157, 8'd158, 8'd78, 8'd155, 8'd103, 8'd127, 8'd90, 8'd119, 8'd165, 8'd145, 8'd83, 8'd123, 8'd162, 8'd167, 8'd162, 8'd176, 8'd110, 8'd149, 8'd86, 8'd168, 8'd111, 8'd68, 8'd65, 8'd67, 8'd161, 8'd165, 8'd156, 8'd113, 8'd129, 8'd145, 8'd126, 8'd136, 8'd85, 8'd93, 8'd93, 8'd126, 8'd166, 8'd77, 8'd165, 8'd93, 8'd112, 8'd170, 8'd174, 8'd137, 8'd130, 8'd120, 8'd166, 8'd180, 8'd141, 8'd126, 8'd114, 8'd162, 8'd155, 8'd123, 8'd108, 8'd144, 8'd128, 8'd96, 8'd164, 8'd71, 8'd101, 8'd171, 8'd123, 8'd84, 8'd156, 8'd123, 8'd106, 8'd104, 8'd192, 8'd111, 8'd130, 8'd152, 8'd140, 8'd120, 8'd143, 8'd119, 8'd162, 8'd122, 8'd72, 8'd148, 8'd83, 8'd80, 8'd91, 8'd156, 8'd70, 8'd78, 8'd86, 8'd87, 8'd87, 8'd93, 8'd80, 8'd94, 8'd143, 8'd80, 8'd137, 8'd125, 8'd127, 8'd179, 8'd121, 8'd137, 8'd214, 8'd146, 8'd183, 8'd107, 8'd122, 8'd164, 8'd154, 8'd114, 8'd138, 8'd99, 8'd112, 8'd139, 8'd78, 8'd143, 8'd119, 8'd93, 8'd86, 8'd125, 8'd106, 8'd122, 8'd142, 8'd142, 8'd131, 8'd152, 8'd156, 8'd158, 8'd185, 8'd191, 8'd176, 8'd122, 8'd136, 8'd141, 8'd133, 8'd101, 8'd63, 8'd127, 8'd58, 8'd90, 8'd117, 8'd100, 8'd83, 8'd162, 8'd162, 8'd94, 8'd127, 8'd94, 8'd78, 8'd84, 8'd62, 8'd93, 8'd140, 8'd75, 8'd65, 8'd67, 8'd77, 8'd177, 8'd88, 8'd93, 8'd106, 8'd119, 8'd97, 8'd75, 8'd80, 8'd55, 8'd102, 8'd90, 8'd68, 8'd144, 8'd72, 8'd116, 8'd154, 8'd139, 8'd132, 8'd114, 8'd108, 8'd138, 8'd114, 8'd122, 8'd95, 8'd56, 8'd121, 8'd95, 8'd136, 8'd154, 8'd157, 8'd121, 8'd69, 8'd84, 8'd113, 8'd67, 8'd83, 8'd146, 8'd59, 8'd92, 8'd63, 8'd116, 8'd70, 8'd151, 8'd213, 8'd189, 8'd119, 8'd165, 8'd74, 8'd79, 8'd132, 8'd48, 8'd80, 8'd74, 8'd64, 8'd55, 8'd83, 8'd58, 8'd146, 8'd121, 8'd85, 8'd83, 8'd104, 8'd125, 8'd106, 8'd75, 8'd61, 8'd143, 8'd115, 8'd71, 8'd115, 8'd99, 8'd149, 8'd176, 8'd95, 8'd101, 8'd86, 8'd113, 8'd82, 8'd110, 8'd72, 8'd82, 8'd94, 8'd93, 8'd137, 8'd129, 8'd76, 8'd67, 8'd67, 8'd134, 8'd92, 8'd148, 8'd155, 8'd134, 8'd124, 8'd65, 8'd149, 8'd75, 8'd83, 8'd95, 8'd172, 8'd128, 8'd142, 8'd147, 8'd72, 8'd111, 8'd134, 8'd140, 8'd115, 8'd114, 8'd91, 8'd92, 8'd117, 8'd152, 8'd97, 8'd116, 8'd154, 8'd120, 8'd80, 8'd123, 8'd72, 8'd68, 8'd136, 8'd75, 8'd133, 8'd69, 8'd158, 8'd153, 8'd154, 8'd151, 8'd157, 8'd92, 8'd123, 8'd120, 8'd159, 8'd127, 8'd84, 8'd99, 8'd129, 8'd102, 8'd116, 8'd134, 8'd155, 8'd113, 8'd74, 8'd147, 8'd72, 8'd126, 8'd153, 8'd89, 8'd71, 8'd90, 8'd172, 8'd76, 8'd130, 8'd108, 8'd142, 8'd134, 8'd120, 8'd169, 8'd91, 8'd176, 8'd114, 8'd88, 8'd111, 8'd180, 8'd103, 8'd141, 8'd142, 8'd109, 8'd145, 8'd177, 8'd108, 8'd152, 8'd104, 8'd150, 8'd158, 8'd142, 8'd93, 8'd110, 8'd146, 8'd146, 8'd146, 8'd142, 8'd106, 8'd170, 8'd135, 8'd97, 8'd104, 8'd100, 8'd156, 8'd147, 8'd147, 8'd116, 8'd76, 8'd102, 8'd156, 8'd176, 8'd101, 8'd133, 8'd133, 8'd168, 8'd118, 8'd147, 8'd91, 8'd107, 8'd84, 8'd65, 8'd164, 8'd157, 8'd116, 8'd81, 8'd97, 8'd132, 8'd98, 8'd133, 8'd165, 8'd187, 8'd158, 8'd166, 8'd167, 8'd131, 8'd117, 8'd158, 8'd184, 8'd165, 8'd115, 8'd174, 8'd114, 8'd103, 8'd163, 8'd158, 8'd161, 8'd169, 8'd121, 8'd151, 8'd75, 8'd123, 8'd111, 8'd117, 8'd106, 8'd98, 8'd160, 8'd163, 8'd119, 8'd117, 8'd162, 8'd172, 8'd148, 8'd102, 8'd141, 8'd148, 8'd163, 8'd84, 8'd122, 8'd131, 8'd148, 8'd154, 8'd91, 8'd154, 8'd76, 8'd82, 8'd125, 8'd118, 8'd100, 8'd165, 8'd92, 8'd132, 8'd78, 8'd141, 8'd94, 8'd103, 8'd151, 8'd160, 8'd132, 8'd141, 8'd75, 8'd78, 8'd101, 8'd114, 8'd79, 8'd80, 8'd115, 8'd110, 8'd70, 8'd94, 8'd113, 8'd128, 8'd132, 8'd100, 8'd162, 8'd133, 8'd110, 8'd106, 8'd71, 8'd153, 8'd150, 8'd94, 8'd80, 8'd165, 8'd139, 8'd165, 8'd106, 8'd84, 8'd74, 8'd160, 8'd155, 8'd77, 8'd87, 8'd67, 8'd122, 8'd88, 8'd103, 8'd82, 8'd100, 8'd151, 8'd106, 8'd113, 8'd138, 8'd130, 8'd135, 8'd135})
) cell_0_0 (
    .clk(clk),
    .input_index(input_index),
    .input_value(input_value),
    .input_result(ground),
    .input_enable(input_enable),
    .output_index(index_0_0_1),
    .output_value(value_0_0_1),
    .output_result(result_0_0_1),
    .output_enable(enable_0_0_1)
);

wire [10-1:0] index_0_1_2;
wire [`DATA_WIDTH-1:0] value_0_1_2;
wire [`DATA_WIDTH*4:0] result_0_1_2;
wire enable_0_1_2;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd84, 8'd71, 8'd118, 8'd166, 8'd155, 8'd113, 8'd100, 8'd137, 8'd94, 8'd59, 8'd115, 8'd133, 8'd150, 8'd73, 8'd59, 8'd74, 8'd108, 8'd118, 8'd127, 8'd79, 8'd139, 8'd76, 8'd129, 8'd138, 8'd111, 8'd106, 8'd107, 8'd170, 8'd134, 8'd89, 8'd81, 8'd122, 8'd130, 8'd148, 8'd88, 8'd129, 8'd138, 8'd132, 8'd169, 8'd122, 8'd129, 8'd167, 8'd101, 8'd149, 8'd164, 8'd161, 8'd156, 8'd100, 8'd183, 8'd173, 8'd120, 8'd165, 8'd151, 8'd122, 8'd78, 8'd160, 8'd125, 8'd78, 8'd149, 8'd123, 8'd125, 8'd159, 8'd124, 8'd97, 8'd124, 8'd149, 8'd153, 8'd82, 8'd112, 8'd117, 8'd80, 8'd114, 8'd98, 8'd78, 8'd78, 8'd117, 8'd129, 8'd128, 8'd97, 8'd128, 8'd112, 8'd151, 8'd160, 8'd110, 8'd146, 8'd127, 8'd84, 8'd146, 8'd151, 8'd102, 8'd111, 8'd113, 8'd99, 8'd99, 8'd82, 8'd154, 8'd139, 8'd118, 8'd136, 8'd168, 8'd142, 8'd84, 8'd165, 8'd79, 8'd116, 8'd102, 8'd65, 8'd138, 8'd77, 8'd106, 8'd110, 8'd77, 8'd158, 8'd75, 8'd160, 8'd126, 8'd138, 8'd126, 8'd133, 8'd128, 8'd95, 8'd143, 8'd125, 8'd118, 8'd99, 8'd112, 8'd125, 8'd117, 8'd164, 8'd106, 8'd84, 8'd164, 8'd93, 8'd77, 8'd111, 8'd111, 8'd98, 8'd132, 8'd169, 8'd131, 8'd146, 8'd60, 8'd171, 8'd180, 8'd121, 8'd133, 8'd157, 8'd135, 8'd101, 8'd107, 8'd87, 8'd139, 8'd96, 8'd98, 8'd107, 8'd174, 8'd162, 8'd158, 8'd119, 8'd119, 8'd104, 8'd167, 8'd75, 8'd151, 8'd62, 8'd91, 8'd143, 8'd71, 8'd102, 8'd132, 8'd109, 8'd175, 8'd170, 8'd163, 8'd161, 8'd74, 8'd132, 8'd133, 8'd80, 8'd125, 8'd69, 8'd84, 8'd104, 8'd97, 8'd61, 8'd154, 8'd122, 8'd75, 8'd116, 8'd146, 8'd86, 8'd96, 8'd109, 8'd144, 8'd161, 8'd115, 8'd148, 8'd101, 8'd148, 8'd167, 8'd128, 8'd153, 8'd160, 8'd155, 8'd143, 8'd137, 8'd103, 8'd86, 8'd145, 8'd88, 8'd67, 8'd98, 8'd59, 8'd99, 8'd77, 8'd149, 8'd108, 8'd157, 8'd152, 8'd121, 8'd43, 8'd101, 8'd81, 8'd100, 8'd147, 8'd133, 8'd162, 8'd88, 8'd115, 8'd163, 8'd73, 8'd85, 8'd91, 8'd115, 8'd93, 8'd114, 8'd88, 8'd69, 8'd112, 8'd95, 8'd149, 8'd129, 8'd80, 8'd162, 8'd140, 8'd120, 8'd71, 8'd144, 8'd44, 8'd137, 8'd105, 8'd123, 8'd87, 8'd162, 8'd109, 8'd85, 8'd120, 8'd94, 8'd126, 8'd106, 8'd151, 8'd90, 8'd63, 8'd108, 8'd97, 8'd91, 8'd122, 8'd134, 8'd178, 8'd93, 8'd93, 8'd89, 8'd168, 8'd148, 8'd101, 8'd149, 8'd121, 8'd126, 8'd124, 8'd164, 8'd160, 8'd144, 8'd109, 8'd140, 8'd61, 8'd78, 8'd68, 8'd89, 8'd96, 8'd116, 8'd106, 8'd111, 8'd164, 8'd114, 8'd88, 8'd165, 8'd105, 8'd170, 8'd180, 8'd109, 8'd126, 8'd83, 8'd119, 8'd158, 8'd128, 8'd106, 8'd98, 8'd71, 8'd166, 8'd95, 8'd141, 8'd91, 8'd65, 8'd55, 8'd98, 8'd71, 8'd110, 8'd82, 8'd143, 8'd84, 8'd83, 8'd79, 8'd137, 8'd70, 8'd167, 8'd142, 8'd158, 8'd154, 8'd109, 8'd122, 8'd85, 8'd173, 8'd109, 8'd86, 8'd135, 8'd88, 8'd82, 8'd166, 8'd125, 8'd122, 8'd122, 8'd125, 8'd137, 8'd109, 8'd76, 8'd95, 8'd80, 8'd125, 8'd106, 8'd124, 8'd63, 8'd88, 8'd147, 8'd134, 8'd93, 8'd172, 8'd136, 8'd132, 8'd101, 8'd147, 8'd71, 8'd123, 8'd111, 8'd118, 8'd84, 8'd124, 8'd148, 8'd151, 8'd74, 8'd134, 8'd113, 8'd153, 8'd168, 8'd145, 8'd139, 8'd102, 8'd147, 8'd98, 8'd114, 8'd151, 8'd136, 8'd67, 8'd94, 8'd173, 8'd127, 8'd101, 8'd89, 8'd118, 8'd97, 8'd99, 8'd111, 8'd64, 8'd99, 8'd174, 8'd105, 8'd140, 8'd154, 8'd121, 8'd108, 8'd150, 8'd185, 8'd99, 8'd137, 8'd97, 8'd119, 8'd144, 8'd141, 8'd68, 8'd116, 8'd87, 8'd169, 8'd128, 8'd98, 8'd139, 8'd176, 8'd94, 8'd88, 8'd108, 8'd77, 8'd150, 8'd156, 8'd113, 8'd95, 8'd107, 8'd188, 8'd131, 8'd160, 8'd119, 8'd141, 8'd100, 8'd115, 8'd113, 8'd59, 8'd92, 8'd120, 8'd129, 8'd94, 8'd138, 8'd166, 8'd167, 8'd170, 8'd149, 8'd136, 8'd121, 8'd93, 8'd50, 8'd104, 8'd114, 8'd111, 8'd82, 8'd69, 8'd105, 8'd136, 8'd113, 8'd124, 8'd122, 8'd118, 8'd120, 8'd110, 8'd143, 8'd62, 8'd129, 8'd152, 8'd147, 8'd109, 8'd136, 8'd114, 8'd129, 8'd104, 8'd89, 8'd158, 8'd142, 8'd105, 8'd103, 8'd101, 8'd111, 8'd82, 8'd119, 8'd114, 8'd56, 8'd138, 8'd165, 8'd167, 8'd99, 8'd132, 8'd139, 8'd96, 8'd132, 8'd110, 8'd69, 8'd80, 8'd131, 8'd129, 8'd130, 8'd139, 8'd106, 8'd93, 8'd174, 8'd171, 8'd134, 8'd79, 8'd103, 8'd92, 8'd68, 8'd155, 8'd144, 8'd120, 8'd141, 8'd168, 8'd148, 8'd163, 8'd106, 8'd173, 8'd184, 8'd149, 8'd106, 8'd142, 8'd122, 8'd134, 8'd109, 8'd91, 8'd170, 8'd124, 8'd140, 8'd104, 8'd174, 8'd99, 8'd140, 8'd127, 8'd126, 8'd59, 8'd112, 8'd77, 8'd69, 8'd86, 8'd126, 8'd128, 8'd120, 8'd175, 8'd149, 8'd151, 8'd126, 8'd125, 8'd149, 8'd110, 8'd160, 8'd170, 8'd140, 8'd155, 8'd121, 8'd106, 8'd107, 8'd135, 8'd148, 8'd140, 8'd90, 8'd134, 8'd117, 8'd93, 8'd162, 8'd69, 8'd91, 8'd93, 8'd83, 8'd111, 8'd95, 8'd98, 8'd157, 8'd84, 8'd90, 8'd121, 8'd115, 8'd120, 8'd133, 8'd147, 8'd95, 8'd158, 8'd131, 8'd82, 8'd114, 8'd101, 8'd121, 8'd112, 8'd151, 8'd119, 8'd95, 8'd138, 8'd97, 8'd102, 8'd106, 8'd82, 8'd45, 8'd144, 8'd92, 8'd126, 8'd157, 8'd131, 8'd103, 8'd176, 8'd167, 8'd122, 8'd151, 8'd178, 8'd117, 8'd85, 8'd91, 8'd159, 8'd121, 8'd98, 8'd98, 8'd115, 8'd110, 8'd147, 8'd133, 8'd137, 8'd86, 8'd99, 8'd95, 8'd118, 8'd45, 8'd126, 8'd90, 8'd142, 8'd76, 8'd142, 8'd147, 8'd146, 8'd133, 8'd85, 8'd162, 8'd98, 8'd118, 8'd75, 8'd127, 8'd125, 8'd150, 8'd105, 8'd95, 8'd44, 8'd143, 8'd98, 8'd149, 8'd126, 8'd112, 8'd113, 8'd94, 8'd140, 8'd46, 8'd63, 8'd60, 8'd60, 8'd92, 8'd48, 8'd55, 8'd66, 8'd99, 8'd76, 8'd62, 8'd60, 8'd136, 8'd124, 8'd61, 8'd66, 8'd105, 8'd68, 8'd131, 8'd97, 8'd100, 8'd97, 8'd158, 8'd117, 8'd125, 8'd157, 8'd98, 8'd114, 8'd103, 8'd78, 8'd134, 8'd44, 8'd27, 8'd72, 8'd112, 8'd26, 8'd93, 8'd39, 8'd106, 8'd42, 8'd95, 8'd108, 8'd59, 8'd151, 8'd135, 8'd97, 8'd77, 8'd157, 8'd93, 8'd142, 8'd68, 8'd79, 8'd161, 8'd135, 8'd106, 8'd153, 8'd93, 8'd78, 8'd130, 8'd64, 8'd67, 8'd40, 8'd37, 8'd43, 8'd50, 8'd123, 8'd91, 8'd46, 8'd75, 8'd68, 8'd47, 8'd117, 8'd88, 8'd146, 8'd123, 8'd127, 8'd82, 8'd110, 8'd117, 8'd110, 8'd170, 8'd76, 8'd103, 8'd122, 8'd100, 8'd116, 8'd115, 8'd64, 8'd138, 8'd68, 8'd146, 8'd83, 8'd139, 8'd71, 8'd131, 8'd118, 8'd159, 8'd110, 8'd103, 8'd111, 8'd92, 8'd118, 8'd120, 8'd68, 8'd98, 8'd111, 8'd141, 8'd75, 8'd133, 8'd147, 8'd118, 8'd164, 8'd115, 8'd140, 8'd142, 8'd126, 8'd100, 8'd164, 8'd128, 8'd137, 8'd91, 8'd95, 8'd136, 8'd133, 8'd107, 8'd91, 8'd110, 8'd125, 8'd120, 8'd149, 8'd88, 8'd154, 8'd128, 8'd155, 8'd90, 8'd104, 8'd93})
) cell_0_1 (
    .clk(clk),
    .input_index(index_0_0_1),
    .input_value(value_0_0_1),
    .input_result(result_0_0_1),
    .input_enable(enable_0_0_1),
    .output_index(index_0_1_2),
    .output_value(value_0_1_2),
    .output_result(result_0_1_2),
    .output_enable(enable_0_1_2)
);

wire [10-1:0] index_0_2_3;
wire [`DATA_WIDTH-1:0] value_0_2_3;
wire [`DATA_WIDTH*4:0] result_0_2_3;
wire enable_0_2_3;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd89, 8'd109, 8'd157, 8'd101, 8'd157, 8'd139, 8'd134, 8'd69, 8'd130, 8'd126, 8'd61, 8'd60, 8'd109, 8'd157, 8'd113, 8'd85, 8'd151, 8'd146, 8'd150, 8'd136, 8'd132, 8'd129, 8'd106, 8'd130, 8'd144, 8'd156, 8'd93, 8'd139, 8'd92, 8'd140, 8'd72, 8'd129, 8'd129, 8'd114, 8'd94, 8'd151, 8'd93, 8'd77, 8'd68, 8'd80, 8'd146, 8'd118, 8'd119, 8'd118, 8'd109, 8'd118, 8'd100, 8'd185, 8'd121, 8'd174, 8'd82, 8'd102, 8'd93, 8'd100, 8'd131, 8'd169, 8'd153, 8'd114, 8'd76, 8'd73, 8'd110, 8'd166, 8'd157, 8'd116, 8'd107, 8'd158, 8'd89, 8'd113, 8'd125, 8'd130, 8'd102, 8'd131, 8'd41, 8'd117, 8'd40, 8'd49, 8'd133, 8'd62, 8'd97, 8'd114, 8'd68, 8'd102, 8'd75, 8'd141, 8'd127, 8'd82, 8'd162, 8'd146, 8'd136, 8'd133, 8'd88, 8'd83, 8'd143, 8'd128, 8'd75, 8'd88, 8'd68, 8'd47, 8'd59, 8'd133, 8'd70, 8'd103, 8'd111, 8'd73, 8'd114, 8'd43, 8'd37, 8'd110, 8'd74, 8'd149, 8'd140, 8'd101, 8'd136, 8'd63, 8'd107, 8'd155, 8'd94, 8'd186, 8'd117, 8'd169, 8'd110, 8'd157, 8'd79, 8'd104, 8'd100, 8'd124, 8'd79, 8'd107, 8'd86, 8'd75, 8'd101, 8'd102, 8'd129, 8'd118, 8'd139, 8'd35, 8'd119, 8'd138, 8'd138, 8'd141, 8'd114, 8'd126, 8'd158, 8'd123, 8'd145, 8'd101, 8'd131, 8'd127, 8'd155, 8'd131, 8'd70, 8'd125, 8'd64, 8'd156, 8'd122, 8'd85, 8'd132, 8'd104, 8'd114, 8'd117, 8'd163, 8'd109, 8'd122, 8'd100, 8'd77, 8'd61, 8'd83, 8'd167, 8'd100, 8'd88, 8'd107, 8'd180, 8'd127, 8'd100, 8'd86, 8'd148, 8'd127, 8'd103, 8'd92, 8'd96, 8'd100, 8'd106, 8'd131, 8'd121, 8'd128, 8'd161, 8'd178, 8'd85, 8'd89, 8'd165, 8'd109, 8'd56, 8'd86, 8'd66, 8'd114, 8'd99, 8'd103, 8'd109, 8'd172, 8'd189, 8'd123, 8'd108, 8'd155, 8'd149, 8'd163, 8'd90, 8'd136, 8'd102, 8'd161, 8'd110, 8'd98, 8'd113, 8'd118, 8'd114, 8'd136, 8'd89, 8'd106, 8'd144, 8'd114, 8'd106, 8'd43, 8'd91, 8'd134, 8'd71, 8'd141, 8'd169, 8'd180, 8'd102, 8'd110, 8'd127, 8'd152, 8'd103, 8'd118, 8'd103, 8'd108, 8'd147, 8'd97, 8'd122, 8'd93, 8'd173, 8'd189, 8'd140, 8'd138, 8'd118, 8'd161, 8'd88, 8'd146, 8'd140, 8'd108, 8'd100, 8'd66, 8'd91, 8'd90, 8'd148, 8'd203, 8'd139, 8'd96, 8'd140, 8'd153, 8'd105, 8'd82, 8'd139, 8'd162, 8'd109, 8'd123, 8'd159, 8'd179, 8'd120, 8'd167, 8'd193, 8'd186, 8'd92, 8'd170, 8'd141, 8'd82, 8'd120, 8'd67, 8'd117, 8'd108, 8'd92, 8'd140, 8'd165, 8'd197, 8'd189, 8'd149, 8'd103, 8'd122, 8'd69, 8'd98, 8'd91, 8'd136, 8'd158, 8'd95, 8'd91, 8'd108, 8'd211, 8'd139, 8'd154, 8'd162, 8'd140, 8'd135, 8'd91, 8'd158, 8'd116, 8'd76, 8'd150, 8'd161, 8'd161, 8'd152, 8'd163, 8'd186, 8'd95, 8'd142, 8'd143, 8'd126, 8'd97, 8'd90, 8'd134, 8'd61, 8'd81, 8'd141, 8'd115, 8'd120, 8'd122, 8'd146, 8'd123, 8'd190, 8'd168, 8'd86, 8'd81, 8'd76, 8'd129, 8'd82, 8'd117, 8'd152, 8'd102, 8'd167, 8'd142, 8'd120, 8'd103, 8'd85, 8'd68, 8'd150, 8'd84, 8'd119, 8'd77, 8'd124, 8'd79, 8'd79, 8'd175, 8'd181, 8'd131, 8'd104, 8'd178, 8'd120, 8'd95, 8'd142, 8'd102, 8'd161, 8'd128, 8'd74, 8'd80, 8'd144, 8'd120, 8'd163, 8'd175, 8'd137, 8'd105, 8'd103, 8'd127, 8'd123, 8'd76, 8'd136, 8'd153, 8'd109, 8'd147, 8'd130, 8'd95, 8'd147, 8'd161, 8'd78, 8'd115, 8'd106, 8'd91, 8'd64, 8'd104, 8'd65, 8'd118, 8'd73, 8'd144, 8'd89, 8'd101, 8'd95, 8'd103, 8'd154, 8'd193, 8'd180, 8'd173, 8'd98, 8'd108, 8'd162, 8'd146, 8'd81, 8'd80, 8'd132, 8'd142, 8'd148, 8'd111, 8'd152, 8'd79, 8'd109, 8'd141, 8'd150, 8'd70, 8'd102, 8'd60, 8'd126, 8'd97, 8'd71, 8'd90, 8'd92, 8'd92, 8'd122, 8'd141, 8'd221, 8'd215, 8'd136, 8'd92, 8'd143, 8'd133, 8'd71, 8'd118, 8'd125, 8'd71, 8'd116, 8'd84, 8'd72, 8'd130, 8'd94, 8'd139, 8'd147, 8'd68, 8'd146, 8'd111, 8'd143, 8'd96, 8'd71, 8'd154, 8'd98, 8'd134, 8'd61, 8'd102, 8'd169, 8'd150, 8'd158, 8'd131, 8'd134, 8'd55, 8'd130, 8'd74, 8'd78, 8'd77, 8'd80, 8'd95, 8'd87, 8'd68, 8'd109, 8'd97, 8'd116, 8'd134, 8'd110, 8'd66, 8'd93, 8'd48, 8'd82, 8'd91, 8'd90, 8'd103, 8'd45, 8'd105, 8'd102, 8'd123, 8'd150, 8'd74, 8'd142, 8'd126, 8'd51, 8'd58, 8'd143, 8'd98, 8'd155, 8'd87, 8'd151, 8'd163, 8'd119, 8'd159, 8'd154, 8'd144, 8'd144, 8'd74, 8'd80, 8'd43, 8'd124, 8'd139, 8'd101, 8'd71, 8'd48, 8'd102, 8'd70, 8'd127, 8'd116, 8'd81, 8'd71, 8'd72, 8'd59, 8'd157, 8'd88, 8'd175, 8'd87, 8'd87, 8'd96, 8'd97, 8'd150, 8'd158, 8'd133, 8'd148, 8'd148, 8'd117, 8'd100, 8'd88, 8'd69, 8'd67, 8'd130, 8'd86, 8'd57, 8'd87, 8'd149, 8'd66, 8'd88, 8'd72, 8'd80, 8'd142, 8'd117, 8'd114, 8'd136, 8'd91, 8'd153, 8'd75, 8'd114, 8'd70, 8'd74, 8'd89, 8'd70, 8'd76, 8'd85, 8'd66, 8'd133, 8'd80, 8'd133, 8'd146, 8'd150, 8'd128, 8'd107, 8'd50, 8'd98, 8'd82, 8'd104, 8'd81, 8'd126, 8'd146, 8'd123, 8'd122, 8'd81, 8'd154, 8'd102, 8'd148, 8'd62, 8'd61, 8'd102, 8'd112, 8'd149, 8'd52, 8'd108, 8'd90, 8'd140, 8'd140, 8'd113, 8'd103, 8'd107, 8'd117, 8'd132, 8'd68, 8'd152, 8'd145, 8'd126, 8'd76, 8'd157, 8'd138, 8'd142, 8'd78, 8'd126, 8'd104, 8'd121, 8'd98, 8'd80, 8'd114, 8'd104, 8'd66, 8'd110, 8'd75, 8'd91, 8'd104, 8'd70, 8'd115, 8'd98, 8'd70, 8'd123, 8'd69, 8'd143, 8'd81, 8'd83, 8'd143, 8'd163, 8'd156, 8'd170, 8'd90, 8'd157, 8'd160, 8'd138, 8'd184, 8'd90, 8'd123, 8'd75, 8'd139, 8'd101, 8'd127, 8'd65, 8'd152, 8'd55, 8'd90, 8'd115, 8'd126, 8'd109, 8'd124, 8'd102, 8'd94, 8'd92, 8'd79, 8'd92, 8'd126, 8'd172, 8'd111, 8'd177, 8'd179, 8'd185, 8'd187, 8'd155, 8'd184, 8'd135, 8'd128, 8'd149, 8'd163, 8'd171, 8'd148, 8'd112, 8'd105, 8'd150, 8'd73, 8'd110, 8'd96, 8'd141, 8'd89, 8'd168, 8'd107, 8'd87, 8'd114, 8'd166, 8'd121, 8'd120, 8'd151, 8'd113, 8'd120, 8'd180, 8'd106, 8'd103, 8'd185, 8'd113, 8'd181, 8'd163, 8'd177, 8'd122, 8'd168, 8'd189, 8'd104, 8'd134, 8'd132, 8'd172, 8'd113, 8'd152, 8'd170, 8'd97, 8'd75, 8'd157, 8'd90, 8'd139, 8'd138, 8'd177, 8'd170, 8'd168, 8'd150, 8'd142, 8'd162, 8'd163, 8'd164, 8'd150, 8'd145, 8'd156, 8'd148, 8'd151, 8'd206, 8'd115, 8'd99, 8'd150, 8'd137, 8'd127, 8'd146, 8'd85, 8'd147, 8'd147, 8'd102, 8'd154, 8'd168, 8'd167, 8'd134, 8'd169, 8'd113, 8'd114, 8'd172, 8'd140, 8'd142, 8'd104, 8'd145, 8'd140, 8'd113, 8'd174, 8'd173, 8'd114, 8'd167, 8'd104, 8'd130, 8'd151, 8'd147, 8'd76, 8'd132, 8'd135, 8'd168, 8'd102, 8'd125, 8'd87, 8'd98, 8'd159, 8'd116, 8'd136, 8'd112, 8'd105, 8'd79, 8'd74, 8'd141, 8'd142, 8'd109, 8'd106, 8'd79, 8'd78, 8'd87, 8'd166, 8'd154, 8'd110, 8'd130, 8'd167, 8'd128, 8'd148, 8'd100, 8'd125, 8'd128})
) cell_0_2 (
    .clk(clk),
    .input_index(index_0_1_2),
    .input_value(value_0_1_2),
    .input_result(result_0_1_2),
    .input_enable(enable_0_1_2),
    .output_index(index_0_2_3),
    .output_value(value_0_2_3),
    .output_result(result_0_2_3),
    .output_enable(enable_0_2_3)
);

wire [10-1:0] index_0_3_4;
wire [`DATA_WIDTH-1:0] value_0_3_4;
wire [`DATA_WIDTH*4:0] result_0_3_4;
wire enable_0_3_4;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd76, 8'd89, 8'd108, 8'd74, 8'd128, 8'd151, 8'd121, 8'd151, 8'd185, 8'd109, 8'd129, 8'd185, 8'd98, 8'd156, 8'd176, 8'd146, 8'd99, 8'd116, 8'd140, 8'd152, 8'd132, 8'd144, 8'd164, 8'd133, 8'd167, 8'd150, 8'd80, 8'd72, 8'd115, 8'd126, 8'd78, 8'd97, 8'd95, 8'd126, 8'd113, 8'd170, 8'd141, 8'd124, 8'd132, 8'd115, 8'd109, 8'd158, 8'd186, 8'd170, 8'd142, 8'd96, 8'd134, 8'd151, 8'd88, 8'd172, 8'd75, 8'd149, 8'd163, 8'd130, 8'd113, 8'd96, 8'd96, 8'd74, 8'd75, 8'd105, 8'd78, 8'd159, 8'd161, 8'd167, 8'd92, 8'd148, 8'd140, 8'd130, 8'd153, 8'd132, 8'd83, 8'd174, 8'd163, 8'd111, 8'd139, 8'd132, 8'd113, 8'd95, 8'd160, 8'd188, 8'd110, 8'd76, 8'd142, 8'd158, 8'd110, 8'd72, 8'd63, 8'd55, 8'd134, 8'd118, 8'd95, 8'd109, 8'd134, 8'd95, 8'd125, 8'd157, 8'd149, 8'd135, 8'd123, 8'd90, 8'd100, 8'd125, 8'd68, 8'd160, 8'd163, 8'd166, 8'd149, 8'd153, 8'd130, 8'd150, 8'd140, 8'd90, 8'd163, 8'd94, 8'd111, 8'd91, 8'd79, 8'd102, 8'd93, 8'd143, 8'd123, 8'd143, 8'd151, 8'd79, 8'd112, 8'd101, 8'd49, 8'd123, 8'd68, 8'd88, 8'd129, 8'd73, 8'd73, 8'd95, 8'd173, 8'd166, 8'd84, 8'd108, 8'd122, 8'd80, 8'd76, 8'd123, 8'd102, 8'd97, 8'd54, 8'd57, 8'd134, 8'd94, 8'd143, 8'd102, 8'd70, 8'd128, 8'd95, 8'd87, 8'd70, 8'd77, 8'd59, 8'd62, 8'd96, 8'd117, 8'd135, 8'd75, 8'd89, 8'd110, 8'd95, 8'd105, 8'd75, 8'd108, 8'd96, 8'd101, 8'd101, 8'd143, 8'd89, 8'd90, 8'd141, 8'd65, 8'd58, 8'd102, 8'd74, 8'd85, 8'd89, 8'd157, 8'd86, 8'd111, 8'd110, 8'd111, 8'd60, 8'd75, 8'd69, 8'd34, 8'd58, 8'd100, 8'd65, 8'd75, 8'd116, 8'd149, 8'd116, 8'd142, 8'd52, 8'd135, 8'd106, 8'd122, 8'd59, 8'd112, 8'd145, 8'd118, 8'd99, 8'd155, 8'd152, 8'd101, 8'd155, 8'd116, 8'd86, 8'd69, 8'd46, 8'd85, 8'd45, 8'd109, 8'd96, 8'd102, 8'd107, 8'd93, 8'd78, 8'd89, 8'd150, 8'd150, 8'd112, 8'd81, 8'd83, 8'd84, 8'd103, 8'd97, 8'd55, 8'd136, 8'd129, 8'd78, 8'd164, 8'd111, 8'd144, 8'd97, 8'd97, 8'd114, 8'd59, 8'd90, 8'd120, 8'd109, 8'd105, 8'd48, 8'd122, 8'd114, 8'd119, 8'd127, 8'd83, 8'd124, 8'd115, 8'd61, 8'd133, 8'd81, 8'd129, 8'd83, 8'd81, 8'd87, 8'd101, 8'd61, 8'd142, 8'd132, 8'd187, 8'd115, 8'd66, 8'd101, 8'd59, 8'd54, 8'd65, 8'd116, 8'd66, 8'd60, 8'd52, 8'd106, 8'd166, 8'd149, 8'd93, 8'd145, 8'd105, 8'd64, 8'd122, 8'd144, 8'd152, 8'd137, 8'd111, 8'd85, 8'd104, 8'd121, 8'd150, 8'd122, 8'd162, 8'd129, 8'd84, 8'd85, 8'd152, 8'd84, 8'd129, 8'd57, 8'd129, 8'd88, 8'd68, 8'd77, 8'd123, 8'd74, 8'd85, 8'd46, 8'd89, 8'd138, 8'd66, 8'd77, 8'd174, 8'd144, 8'd116, 8'd158, 8'd144, 8'd139, 8'd127, 8'd161, 8'd144, 8'd115, 8'd96, 8'd146, 8'd144, 8'd77, 8'd95, 8'd146, 8'd73, 8'd89, 8'd134, 8'd78, 8'd176, 8'd169, 8'd88, 8'd132, 8'd41, 8'd112, 8'd110, 8'd174, 8'd120, 8'd138, 8'd119, 8'd148, 8'd190, 8'd111, 8'd109, 8'd157, 8'd92, 8'd120, 8'd153, 8'd130, 8'd158, 8'd83, 8'd124, 8'd91, 8'd178, 8'd118, 8'd130, 8'd178, 8'd90, 8'd143, 8'd70, 8'd48, 8'd91, 8'd74, 8'd170, 8'd92, 8'd96, 8'd168, 8'd116, 8'd162, 8'd156, 8'd144, 8'd152, 8'd133, 8'd121, 8'd42, 8'd85, 8'd112, 8'd90, 8'd133, 8'd173, 8'd109, 8'd147, 8'd166, 8'd117, 8'd93, 8'd173, 8'd99, 8'd121, 8'd137, 8'd85, 8'd72, 8'd70, 8'd132, 8'd87, 8'd99, 8'd151, 8'd129, 8'd174, 8'd153, 8'd102, 8'd106, 8'd41, 8'd117, 8'd157, 8'd131, 8'd103, 8'd107, 8'd135, 8'd207, 8'd128, 8'd176, 8'd101, 8'd160, 8'd99, 8'd174, 8'd130, 8'd48, 8'd65, 8'd134, 8'd56, 8'd143, 8'd94, 8'd136, 8'd155, 8'd114, 8'd127, 8'd163, 8'd107, 8'd167, 8'd109, 8'd148, 8'd94, 8'd123, 8'd184, 8'd166, 8'd149, 8'd100, 8'd142, 8'd120, 8'd187, 8'd194, 8'd89, 8'd120, 8'd104, 8'd113, 8'd42, 8'd107, 8'd99, 8'd99, 8'd85, 8'd116, 8'd106, 8'd102, 8'd180, 8'd145, 8'd159, 8'd168, 8'd127, 8'd124, 8'd150, 8'd115, 8'd129, 8'd179, 8'd182, 8'd78, 8'd138, 8'd173, 8'd155, 8'd117, 8'd89, 8'd137, 8'd86, 8'd112, 8'd125, 8'd118, 8'd111, 8'd112, 8'd155, 8'd142, 8'd67, 8'd150, 8'd131, 8'd126, 8'd126, 8'd78, 8'd150, 8'd173, 8'd86, 8'd172, 8'd165, 8'd136, 8'd129, 8'd127, 8'd158, 8'd125, 8'd131, 8'd177, 8'd91, 8'd104, 8'd98, 8'd97, 8'd47, 8'd45, 8'd134, 8'd153, 8'd89, 8'd135, 8'd107, 8'd71, 8'd108, 8'd80, 8'd121, 8'd67, 8'd165, 8'd141, 8'd113, 8'd119, 8'd69, 8'd107, 8'd68, 8'd94, 8'd95, 8'd161, 8'd91, 8'd135, 8'd182, 8'd109, 8'd123, 8'd83, 8'd83, 8'd76, 8'd137, 8'd135, 8'd154, 8'd68, 8'd139, 8'd104, 8'd138, 8'd146, 8'd86, 8'd60, 8'd129, 8'd106, 8'd154, 8'd71, 8'd90, 8'd117, 8'd111, 8'd105, 8'd86, 8'd73, 8'd164, 8'd114, 8'd144, 8'd134, 8'd89, 8'd116, 8'd77, 8'd134, 8'd139, 8'd107, 8'd66, 8'd161, 8'd104, 8'd114, 8'd78, 8'd87, 8'd67, 8'd50, 8'd153, 8'd104, 8'd80, 8'd126, 8'd143, 8'd105, 8'd116, 8'd73, 8'd166, 8'd77, 8'd173, 8'd101, 8'd149, 8'd145, 8'd108, 8'd155, 8'd94, 8'd166, 8'd93, 8'd123, 8'd151, 8'd158, 8'd64, 8'd58, 8'd74, 8'd65, 8'd47, 8'd55, 8'd96, 8'd83, 8'd83, 8'd134, 8'd132, 8'd78, 8'd107, 8'd172, 8'd98, 8'd115, 8'd173, 8'd174, 8'd128, 8'd156, 8'd134, 8'd104, 8'd101, 8'd129, 8'd209, 8'd146, 8'd106, 8'd109, 8'd146, 8'd134, 8'd105, 8'd101, 8'd85, 8'd50, 8'd124, 8'd60, 8'd128, 8'd90, 8'd77, 8'd68, 8'd112, 8'd129, 8'd157, 8'd122, 8'd85, 8'd111, 8'd115, 8'd168, 8'd96, 8'd145, 8'd89, 8'd120, 8'd154, 8'd164, 8'd194, 8'd188, 8'd165, 8'd144, 8'd66, 8'd114, 8'd70, 8'd106, 8'd126, 8'd103, 8'd81, 8'd44, 8'd95, 8'd59, 8'd65, 8'd68, 8'd112, 8'd100, 8'd156, 8'd150, 8'd83, 8'd106, 8'd132, 8'd114, 8'd171, 8'd189, 8'd154, 8'd118, 8'd125, 8'd116, 8'd126, 8'd134, 8'd87, 8'd115, 8'd111, 8'd115, 8'd49, 8'd62, 8'd114, 8'd44, 8'd114, 8'd128, 8'd157, 8'd148, 8'd92, 8'd155, 8'd80, 8'd107, 8'd144, 8'd119, 8'd125, 8'd118, 8'd71, 8'd151, 8'd162, 8'd97, 8'd97, 8'd151, 8'd134, 8'd168, 8'd93, 8'd136, 8'd160, 8'd175, 8'd155, 8'd62, 8'd91, 8'd150, 8'd122, 8'd151, 8'd97, 8'd120, 8'd163, 8'd153, 8'd122, 8'd133, 8'd98, 8'd142, 8'd157, 8'd80, 8'd113, 8'd90, 8'd62, 8'd152, 8'd79, 8'd68, 8'd110, 8'd153, 8'd110, 8'd119, 8'd103, 8'd101, 8'd97, 8'd97, 8'd64, 8'd105, 8'd152, 8'd123, 8'd115, 8'd59, 8'd126, 8'd76, 8'd117, 8'd97, 8'd108, 8'd116, 8'd105, 8'd80, 8'd166, 8'd102, 8'd100, 8'd169, 8'd159, 8'd111, 8'd76, 8'd159, 8'd112, 8'd114, 8'd76, 8'd101, 8'd142, 8'd140, 8'd97, 8'd87, 8'd115, 8'd77, 8'd168, 8'd148, 8'd74, 8'd162, 8'd149, 8'd134, 8'd114, 8'd114})
) cell_0_3 (
    .clk(clk),
    .input_index(index_0_2_3),
    .input_value(value_0_2_3),
    .input_result(result_0_2_3),
    .input_enable(enable_0_2_3),
    .output_index(index_0_3_4),
    .output_value(value_0_3_4),
    .output_result(result_0_3_4),
    .output_enable(enable_0_3_4)
);

wire [10-1:0] index_0_4_5;
wire [`DATA_WIDTH-1:0] value_0_4_5;
wire [`DATA_WIDTH*4:0] result_0_4_5;
wire enable_0_4_5;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd80, 8'd161, 8'd76, 8'd86, 8'd113, 8'd89, 8'd110, 8'd84, 8'd117, 8'd142, 8'd97, 8'd73, 8'd48, 8'd139, 8'd65, 8'd140, 8'd132, 8'd99, 8'd121, 8'd67, 8'd83, 8'd133, 8'd141, 8'd161, 8'd129, 8'd144, 8'd100, 8'd167, 8'd73, 8'd123, 8'd93, 8'd94, 8'd83, 8'd91, 8'd99, 8'd91, 8'd110, 8'd144, 8'd90, 8'd154, 8'd134, 8'd74, 8'd77, 8'd157, 8'd76, 8'd142, 8'd119, 8'd93, 8'd118, 8'd129, 8'd136, 8'd116, 8'd153, 8'd72, 8'd108, 8'd135, 8'd137, 8'd76, 8'd153, 8'd108, 8'd100, 8'd130, 8'd92, 8'd98, 8'd117, 8'd115, 8'd111, 8'd155, 8'd188, 8'd190, 8'd160, 8'd189, 8'd203, 8'd137, 8'd175, 8'd159, 8'd181, 8'd102, 8'd171, 8'd102, 8'd161, 8'd154, 8'd164, 8'd156, 8'd168, 8'd101, 8'd120, 8'd117, 8'd102, 8'd118, 8'd124, 8'd147, 8'd118, 8'd118, 8'd138, 8'd82, 8'd151, 8'd146, 8'd156, 8'd132, 8'd153, 8'd171, 8'd134, 8'd114, 8'd136, 8'd156, 8'd173, 8'd127, 8'd130, 8'd119, 8'd82, 8'd160, 8'd109, 8'd97, 8'd142, 8'd109, 8'd67, 8'd150, 8'd107, 8'd112, 8'd132, 8'd87, 8'd102, 8'd109, 8'd145, 8'd102, 8'd117, 8'd91, 8'd96, 8'd114, 8'd117, 8'd80, 8'd113, 8'd178, 8'd134, 8'd194, 8'd198, 8'd137, 8'd100, 8'd135, 8'd102, 8'd142, 8'd163, 8'd135, 8'd146, 8'd110, 8'd155, 8'd165, 8'd107, 8'd110, 8'd118, 8'd134, 8'd125, 8'd116, 8'd140, 8'd80, 8'd118, 8'd128, 8'd104, 8'd149, 8'd92, 8'd94, 8'd94, 8'd101, 8'd105, 8'd102, 8'd110, 8'd167, 8'd101, 8'd162, 8'd104, 8'd151, 8'd66, 8'd74, 8'd94, 8'd96, 8'd144, 8'd106, 8'd162, 8'd181, 8'd159, 8'd162, 8'd107, 8'd125, 8'd158, 8'd150, 8'd77, 8'd147, 8'd78, 8'd73, 8'd169, 8'd156, 8'd110, 8'd93, 8'd162, 8'd117, 8'd148, 8'd143, 8'd90, 8'd91, 8'd105, 8'd160, 8'd156, 8'd181, 8'd173, 8'd153, 8'd163, 8'd95, 8'd168, 8'd96, 8'd156, 8'd81, 8'd124, 8'd139, 8'd114, 8'd115, 8'd144, 8'd147, 8'd172, 8'd175, 8'd147, 8'd134, 8'd104, 8'd96, 8'd133, 8'd87, 8'd122, 8'd75, 8'd127, 8'd103, 8'd117, 8'd133, 8'd151, 8'd131, 8'd172, 8'd133, 8'd139, 8'd150, 8'd108, 8'd60, 8'd66, 8'd124, 8'd102, 8'd71, 8'd134, 8'd102, 8'd124, 8'd159, 8'd137, 8'd163, 8'd85, 8'd95, 8'd76, 8'd110, 8'd91, 8'd116, 8'd126, 8'd124, 8'd138, 8'd126, 8'd110, 8'd138, 8'd138, 8'd134, 8'd136, 8'd135, 8'd139, 8'd64, 8'd79, 8'd104, 8'd88, 8'd89, 8'd129, 8'd115, 8'd143, 8'd187, 8'd108, 8'd151, 8'd127, 8'd116, 8'd107, 8'd100, 8'd77, 8'd116, 8'd175, 8'd83, 8'd113, 8'd100, 8'd151, 8'd123, 8'd111, 8'd154, 8'd81, 8'd57, 8'd45, 8'd123, 8'd127, 8'd44, 8'd62, 8'd110, 8'd59, 8'd99, 8'd162, 8'd134, 8'd169, 8'd94, 8'd124, 8'd73, 8'd129, 8'd30, 8'd119, 8'd113, 8'd123, 8'd103, 8'd166, 8'd158, 8'd123, 8'd105, 8'd123, 8'd84, 8'd136, 8'd112, 8'd101, 8'd77, 8'd66, 8'd81, 8'd57, 8'd39, 8'd58, 8'd107, 8'd147, 8'd100, 8'd156, 8'd108, 8'd118, 8'd73, 8'd56, 8'd72, 8'd104, 8'd99, 8'd160, 8'd178, 8'd112, 8'd104, 8'd167, 8'd151, 8'd65, 8'd125, 8'd114, 8'd141, 8'd127, 8'd126, 8'd163, 8'd147, 8'd150, 8'd54, 8'd47, 8'd146, 8'd93, 8'd96, 8'd94, 8'd120, 8'd83, 8'd163, 8'd97, 8'd77, 8'd122, 8'd59, 8'd77, 8'd132, 8'd116, 8'd99, 8'd160, 8'd70, 8'd123, 8'd182, 8'd101, 8'd188, 8'd135, 8'd110, 8'd113, 8'd113, 8'd108, 8'd73, 8'd68, 8'd127, 8'd148, 8'd158, 8'd148, 8'd87, 8'd130, 8'd110, 8'd124, 8'd118, 8'd118, 8'd38, 8'd83, 8'd118, 8'd45, 8'd92, 8'd123, 8'd102, 8'd120, 8'd109, 8'd135, 8'd197, 8'd128, 8'd160, 8'd162, 8'd174, 8'd106, 8'd120, 8'd130, 8'd151, 8'd142, 8'd96, 8'd162, 8'd139, 8'd117, 8'd146, 8'd100, 8'd92, 8'd69, 8'd77, 8'd94, 8'd59, 8'd61, 8'd43, 8'd71, 8'd78, 8'd162, 8'd136, 8'd165, 8'd187, 8'd142, 8'd134, 8'd147, 8'd135, 8'd107, 8'd146, 8'd121, 8'd94, 8'd120, 8'd87, 8'd110, 8'd98, 8'd73, 8'd154, 8'd144, 8'd106, 8'd187, 8'd168, 8'd140, 8'd53, 8'd68, 8'd96, 8'd112, 8'd81, 8'd110, 8'd114, 8'd150, 8'd128, 8'd159, 8'd128, 8'd96, 8'd115, 8'd89, 8'd77, 8'd66, 8'd124, 8'd142, 8'd93, 8'd166, 8'd141, 8'd70, 8'd82, 8'd159, 8'd150, 8'd169, 8'd167, 8'd97, 8'd150, 8'd57, 8'd84, 8'd52, 8'd100, 8'd133, 8'd113, 8'd85, 8'd169, 8'd156, 8'd140, 8'd98, 8'd116, 8'd146, 8'd106, 8'd103, 8'd79, 8'd103, 8'd121, 8'd134, 8'd137, 8'd82, 8'd97, 8'd94, 8'd153, 8'd161, 8'd179, 8'd73, 8'd76, 8'd119, 8'd147, 8'd48, 8'd130, 8'd72, 8'd136, 8'd89, 8'd168, 8'd70, 8'd91, 8'd106, 8'd66, 8'd136, 8'd128, 8'd156, 8'd106, 8'd140, 8'd108, 8'd143, 8'd129, 8'd72, 8'd158, 8'd77, 8'd137, 8'd188, 8'd149, 8'd83, 8'd136, 8'd88, 8'd68, 8'd64, 8'd134, 8'd70, 8'd167, 8'd134, 8'd163, 8'd99, 8'd107, 8'd118, 8'd67, 8'd108, 8'd151, 8'd123, 8'd109, 8'd128, 8'd131, 8'd136, 8'd73, 8'd116, 8'd101, 8'd161, 8'd122, 8'd188, 8'd162, 8'd72, 8'd102, 8'd151, 8'd156, 8'd128, 8'd86, 8'd110, 8'd185, 8'd164, 8'd108, 8'd152, 8'd147, 8'd108, 8'd115, 8'd91, 8'd75, 8'd106, 8'd105, 8'd88, 8'd108, 8'd129, 8'd129, 8'd164, 8'd150, 8'd178, 8'd173, 8'd172, 8'd190, 8'd136, 8'd99, 8'd153, 8'd112, 8'd96, 8'd96, 8'd87, 8'd137, 8'd87, 8'd107, 8'd124, 8'd87, 8'd85, 8'd147, 8'd146, 8'd127, 8'd98, 8'd86, 8'd74, 8'd155, 8'd118, 8'd163, 8'd162, 8'd90, 8'd110, 8'd89, 8'd109, 8'd168, 8'd86, 8'd148, 8'd163, 8'd150, 8'd81, 8'd112, 8'd131, 8'd127, 8'd147, 8'd142, 8'd151, 8'd101, 8'd93, 8'd117, 8'd166, 8'd122, 8'd100, 8'd151, 8'd145, 8'd147, 8'd161, 8'd134, 8'd160, 8'd119, 8'd142, 8'd79, 8'd99, 8'd171, 8'd112, 8'd173, 8'd182, 8'd157, 8'd93, 8'd156, 8'd94, 8'd70, 8'd102, 8'd131, 8'd108, 8'd103, 8'd163, 8'd150, 8'd107, 8'd84, 8'd115, 8'd135, 8'd95, 8'd174, 8'd85, 8'd172, 8'd169, 8'd108, 8'd88, 8'd107, 8'd114, 8'd124, 8'd141, 8'd125, 8'd151, 8'd117, 8'd128, 8'd196, 8'd172, 8'd177, 8'd197, 8'd101, 8'd100, 8'd93, 8'd171, 8'd171, 8'd129, 8'd176, 8'd179, 8'd105, 8'd101, 8'd133, 8'd93, 8'd93, 8'd157, 8'd94, 8'd130, 8'd92, 8'd92, 8'd81, 8'd110, 8'd188, 8'd109, 8'd167, 8'd112, 8'd114, 8'd118, 8'd131, 8'd111, 8'd110, 8'd149, 8'd121, 8'd116, 8'd150, 8'd130, 8'd157, 8'd146, 8'd126, 8'd150, 8'd139, 8'd90, 8'd154, 8'd93, 8'd151, 8'd141, 8'd86, 8'd79, 8'd81, 8'd99, 8'd124, 8'd99, 8'd159, 8'd117, 8'd165, 8'd81, 8'd91, 8'd87, 8'd102, 8'd143, 8'd110, 8'd97, 8'd113, 8'd141, 8'd163, 8'd154, 8'd134, 8'd144, 8'd80, 8'd120, 8'd155, 8'd135, 8'd84, 8'd146, 8'd166, 8'd155, 8'd100, 8'd80, 8'd105, 8'd90, 8'd124, 8'd108, 8'd72, 8'd78, 8'd116, 8'd149, 8'd105, 8'd156, 8'd139, 8'd109, 8'd157, 8'd147, 8'd105, 8'd129, 8'd103, 8'd88, 8'd96, 8'd71, 8'd128, 8'd146, 8'd122})
) cell_0_4 (
    .clk(clk),
    .input_index(index_0_3_4),
    .input_value(value_0_3_4),
    .input_result(result_0_3_4),
    .input_enable(enable_0_3_4),
    .output_index(index_0_4_5),
    .output_value(value_0_4_5),
    .output_result(result_0_4_5),
    .output_enable(enable_0_4_5)
);

wire [10-1:0] index_0_5_6;
wire [`DATA_WIDTH-1:0] value_0_5_6;
wire [`DATA_WIDTH*4:0] result_0_5_6;
wire enable_0_5_6;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd84, 8'd90, 8'd146, 8'd111, 8'd63, 8'd97, 8'd111, 8'd98, 8'd74, 8'd64, 8'd121, 8'd140, 8'd150, 8'd143, 8'd144, 8'd97, 8'd65, 8'd71, 8'd98, 8'd105, 8'd92, 8'd101, 8'd104, 8'd163, 8'd128, 8'd81, 8'd95, 8'd136, 8'd89, 8'd85, 8'd123, 8'd143, 8'd122, 8'd74, 8'd130, 8'd120, 8'd74, 8'd109, 8'd59, 8'd103, 8'd125, 8'd119, 8'd75, 8'd67, 8'd68, 8'd94, 8'd89, 8'd131, 8'd126, 8'd133, 8'd132, 8'd64, 8'd70, 8'd103, 8'd118, 8'd142, 8'd92, 8'd154, 8'd89, 8'd160, 8'd152, 8'd130, 8'd95, 8'd106, 8'd145, 8'd90, 8'd100, 8'd120, 8'd128, 8'd59, 8'd67, 8'd110, 8'd93, 8'd54, 8'd133, 8'd102, 8'd90, 8'd62, 8'd113, 8'd136, 8'd96, 8'd122, 8'd162, 8'd132, 8'd130, 8'd112, 8'd112, 8'd138, 8'd151, 8'd138, 8'd129, 8'd147, 8'd82, 8'd77, 8'd77, 8'd111, 8'd90, 8'd114, 8'd108, 8'd83, 8'd94, 8'd143, 8'd160, 8'd101, 8'd46, 8'd74, 8'd58, 8'd51, 8'd131, 8'd111, 8'd144, 8'd153, 8'd112, 8'd92, 8'd111, 8'd68, 8'd69, 8'd94, 8'd69, 8'd109, 8'd127, 8'd104, 8'd153, 8'd84, 8'd143, 8'd101, 8'd116, 8'd135, 8'd103, 8'd131, 8'd124, 8'd109, 8'd106, 8'd149, 8'd148, 8'd149, 8'd139, 8'd104, 8'd104, 8'd144, 8'd125, 8'd137, 8'd90, 8'd128, 8'd144, 8'd128, 8'd85, 8'd79, 8'd105, 8'd89, 8'd135, 8'd113, 8'd135, 8'd176, 8'd101, 8'd81, 8'd107, 8'd138, 8'd107, 8'd156, 8'd135, 8'd87, 8'd108, 8'd132, 8'd159, 8'd128, 8'd99, 8'd173, 8'd86, 8'd88, 8'd67, 8'd63, 8'd110, 8'd143, 8'd91, 8'd122, 8'd95, 8'd161, 8'd119, 8'd171, 8'd124, 8'd129, 8'd149, 8'd87, 8'd154, 8'd132, 8'd83, 8'd145, 8'd106, 8'd127, 8'd165, 8'd154, 8'd140, 8'd117, 8'd112, 8'd98, 8'd157, 8'd105, 8'd120, 8'd92, 8'd114, 8'd91, 8'd105, 8'd97, 8'd80, 8'd86, 8'd129, 8'd148, 8'd150, 8'd93, 8'd101, 8'd185, 8'd139, 8'd172, 8'd157, 8'd160, 8'd149, 8'd138, 8'd156, 8'd70, 8'd120, 8'd127, 8'd131, 8'd113, 8'd156, 8'd123, 8'd96, 8'd60, 8'd91, 8'd135, 8'd138, 8'd165, 8'd97, 8'd146, 8'd117, 8'd108, 8'd80, 8'd128, 8'd153, 8'd107, 8'd97, 8'd107, 8'd158, 8'd185, 8'd99, 8'd100, 8'd91, 8'd97, 8'd71, 8'd95, 8'd159, 8'd165, 8'd159, 8'd66, 8'd125, 8'd148, 8'd164, 8'd123, 8'd88, 8'd127, 8'd76, 8'd143, 8'd117, 8'd122, 8'd158, 8'd152, 8'd123, 8'd116, 8'd125, 8'd143, 8'd95, 8'd138, 8'd94, 8'd148, 8'd66, 8'd119, 8'd152, 8'd178, 8'd150, 8'd107, 8'd132, 8'd147, 8'd120, 8'd95, 8'd97, 8'd98, 8'd72, 8'd126, 8'd151, 8'd69, 8'd131, 8'd74, 8'd85, 8'd82, 8'd129, 8'd181, 8'd151, 8'd171, 8'd130, 8'd116, 8'd98, 8'd63, 8'd117, 8'd105, 8'd114, 8'd100, 8'd148, 8'd84, 8'd120, 8'd110, 8'd118, 8'd120, 8'd77, 8'd113, 8'd87, 8'd135, 8'd84, 8'd102, 8'd71, 8'd56, 8'd121, 8'd161, 8'd148, 8'd111, 8'd153, 8'd132, 8'd89, 8'd94, 8'd102, 8'd87, 8'd133, 8'd106, 8'd146, 8'd113, 8'd169, 8'd100, 8'd111, 8'd75, 8'd98, 8'd109, 8'd126, 8'd76, 8'd127, 8'd56, 8'd49, 8'd135, 8'd106, 8'd139, 8'd123, 8'd170, 8'd189, 8'd96, 8'd120, 8'd109, 8'd93, 8'd103, 8'd130, 8'd70, 8'd144, 8'd61, 8'd87, 8'd132, 8'd146, 8'd157, 8'd157, 8'd117, 8'd106, 8'd175, 8'd114, 8'd75, 8'd72, 8'd125, 8'd144, 8'd74, 8'd148, 8'd102, 8'd130, 8'd192, 8'd105, 8'd133, 8'd91, 8'd122, 8'd64, 8'd66, 8'd62, 8'd52, 8'd70, 8'd39, 8'd136, 8'd152, 8'd139, 8'd79, 8'd121, 8'd87, 8'd151, 8'd138, 8'd191, 8'd128, 8'd84, 8'd112, 8'd73, 8'd114, 8'd105, 8'd88, 8'd113, 8'd164, 8'd127, 8'd191, 8'd73, 8'd126, 8'd137, 8'd144, 8'd106, 8'd81, 8'd78, 8'd58, 8'd90, 8'd104, 8'd161, 8'd162, 8'd147, 8'd121, 8'd92, 8'd172, 8'd163, 8'd188, 8'd88, 8'd148, 8'd150, 8'd61, 8'd87, 8'd64, 8'd87, 8'd152, 8'd159, 8'd113, 8'd103, 8'd90, 8'd97, 8'd115, 8'd98, 8'd110, 8'd126, 8'd121, 8'd88, 8'd166, 8'd105, 8'd150, 8'd100, 8'd95, 8'd148, 8'd178, 8'd154, 8'd102, 8'd171, 8'd154, 8'd155, 8'd119, 8'd123, 8'd72, 8'd98, 8'd192, 8'd140, 8'd146, 8'd136, 8'd161, 8'd170, 8'd179, 8'd157, 8'd105, 8'd85, 8'd133, 8'd71, 8'd79, 8'd154, 8'd117, 8'd139, 8'd142, 8'd108, 8'd93, 8'd148, 8'd148, 8'd98, 8'd167, 8'd138, 8'd90, 8'd122, 8'd130, 8'd95, 8'd152, 8'd126, 8'd168, 8'd158, 8'd99, 8'd155, 8'd134, 8'd93, 8'd105, 8'd103, 8'd154, 8'd166, 8'd123, 8'd96, 8'd91, 8'd104, 8'd142, 8'd137, 8'd155, 8'd174, 8'd132, 8'd108, 8'd125, 8'd141, 8'd99, 8'd70, 8'd120, 8'd93, 8'd77, 8'd115, 8'd111, 8'd114, 8'd134, 8'd139, 8'd109, 8'd167, 8'd175, 8'd126, 8'd96, 8'd127, 8'd131, 8'd111, 8'd146, 8'd148, 8'd163, 8'd150, 8'd158, 8'd165, 8'd109, 8'd130, 8'd106, 8'd114, 8'd87, 8'd73, 8'd129, 8'd77, 8'd107, 8'd67, 8'd91, 8'd66, 8'd82, 8'd132, 8'd124, 8'd155, 8'd81, 8'd130, 8'd144, 8'd150, 8'd125, 8'd137, 8'd98, 8'd91, 8'd100, 8'd95, 8'd99, 8'd149, 8'd110, 8'd98, 8'd118, 8'd130, 8'd88, 8'd85, 8'd147, 8'd97, 8'd130, 8'd132, 8'd91, 8'd132, 8'd134, 8'd99, 8'd122, 8'd172, 8'd153, 8'd102, 8'd112, 8'd108, 8'd58, 8'd99, 8'd167, 8'd155, 8'd132, 8'd120, 8'd92, 8'd136, 8'd170, 8'd90, 8'd141, 8'd163, 8'd144, 8'd78, 8'd143, 8'd103, 8'd133, 8'd160, 8'd95, 8'd160, 8'd121, 8'd155, 8'd141, 8'd164, 8'd77, 8'd88, 8'd145, 8'd126, 8'd140, 8'd157, 8'd70, 8'd152, 8'd147, 8'd161, 8'd145, 8'd84, 8'd124, 8'd132, 8'd128, 8'd165, 8'd170, 8'd113, 8'd168, 8'd133, 8'd166, 8'd87, 8'd89, 8'd158, 8'd133, 8'd106, 8'd130, 8'd152, 8'd152, 8'd77, 8'd111, 8'd138, 8'd157, 8'd104, 8'd110, 8'd104, 8'd130, 8'd87, 8'd102, 8'd104, 8'd121, 8'd139, 8'd134, 8'd143, 8'd145, 8'd135, 8'd113, 8'd147, 8'd169, 8'd178, 8'd106, 8'd175, 8'd111, 8'd111, 8'd106, 8'd93, 8'd167, 8'd145, 8'd124, 8'd169, 8'd105, 8'd161, 8'd73, 8'd147, 8'd116, 8'd66, 8'd136, 8'd138, 8'd142, 8'd105, 8'd119, 8'd146, 8'd111, 8'd100, 8'd107, 8'd160, 8'd142, 8'd139, 8'd171, 8'd164, 8'd177, 8'd160, 8'd119, 8'd129, 8'd145, 8'd128, 8'd104, 8'd153, 8'd89, 8'd139, 8'd101, 8'd145, 8'd115, 8'd107, 8'd168, 8'd187, 8'd94, 8'd116, 8'd118, 8'd137, 8'd167, 8'd109, 8'd132, 8'd131, 8'd164, 8'd137, 8'd119, 8'd117, 8'd184, 8'd97, 8'd131, 8'd135, 8'd129, 8'd100, 8'd119, 8'd111, 8'd80, 8'd120, 8'd85, 8'd86, 8'd136, 8'd138, 8'd168, 8'd83, 8'd179, 8'd105, 8'd133, 8'd105, 8'd171, 8'd105, 8'd158, 8'd144, 8'd92, 8'd125, 8'd162, 8'd163, 8'd99, 8'd113, 8'd131, 8'd173, 8'd97, 8'd132, 8'd87, 8'd117, 8'd152, 8'd90, 8'd86, 8'd125, 8'd135, 8'd110, 8'd82, 8'd157, 8'd96, 8'd153, 8'd137, 8'd108, 8'd77, 8'd85, 8'd170, 8'd142, 8'd165, 8'd124, 8'd98, 8'd160, 8'd80, 8'd95, 8'd139, 8'd114, 8'd159, 8'd83, 8'd71, 8'd121, 8'd144, 8'd75, 8'd166})
) cell_0_5 (
    .clk(clk),
    .input_index(index_0_4_5),
    .input_value(value_0_4_5),
    .input_result(result_0_4_5),
    .input_enable(enable_0_4_5),
    .output_index(index_0_5_6),
    .output_value(value_0_5_6),
    .output_result(result_0_5_6),
    .output_enable(enable_0_5_6)
);

wire [10-1:0] index_0_6_7;
wire [`DATA_WIDTH-1:0] value_0_6_7;
wire [`DATA_WIDTH*4:0] result_0_6_7;
wire enable_0_6_7;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd108, 8'd163, 8'd139, 8'd117, 8'd163, 8'd123, 8'd139, 8'd138, 8'd110, 8'd106, 8'd130, 8'd83, 8'd135, 8'd94, 8'd126, 8'd147, 8'd142, 8'd96, 8'd117, 8'd88, 8'd99, 8'd124, 8'd126, 8'd162, 8'd137, 8'd124, 8'd93, 8'd106, 8'd122, 8'd125, 8'd118, 8'd129, 8'd154, 8'd142, 8'd105, 8'd110, 8'd98, 8'd104, 8'd193, 8'd140, 8'd122, 8'd119, 8'd183, 8'd136, 8'd126, 8'd122, 8'd187, 8'd136, 8'd140, 8'd163, 8'd122, 8'd105, 8'd119, 8'd136, 8'd88, 8'd106, 8'd155, 8'd96, 8'd152, 8'd104, 8'd161, 8'd115, 8'd99, 8'd162, 8'd143, 8'd156, 8'd124, 8'd121, 8'd150, 8'd162, 8'd94, 8'd135, 8'd122, 8'd174, 8'd86, 8'd142, 8'd80, 8'd140, 8'd73, 8'd120, 8'd78, 8'd156, 8'd73, 8'd141, 8'd163, 8'd103, 8'd120, 8'd145, 8'd80, 8'd100, 8'd98, 8'd121, 8'd168, 8'd89, 8'd98, 8'd98, 8'd137, 8'd155, 8'd84, 8'd135, 8'd172, 8'd130, 8'd115, 8'd130, 8'd120, 8'd180, 8'd149, 8'd143, 8'd164, 8'd164, 8'd162, 8'd137, 8'd127, 8'd75, 8'd136, 8'd123, 8'd89, 8'd140, 8'd99, 8'd143, 8'd107, 8'd117, 8'd79, 8'd108, 8'd80, 8'd99, 8'd156, 8'd91, 8'd127, 8'd156, 8'd159, 8'd141, 8'd99, 8'd165, 8'd80, 8'd144, 8'd139, 8'd161, 8'd92, 8'd77, 8'd122, 8'd154, 8'd92, 8'd108, 8'd70, 8'd81, 8'd152, 8'd156, 8'd159, 8'd136, 8'd74, 8'd101, 8'd112, 8'd77, 8'd108, 8'd104, 8'd113, 8'd79, 8'd122, 8'd171, 8'd113, 8'd98, 8'd149, 8'd119, 8'd101, 8'd86, 8'd77, 8'd102, 8'd154, 8'd126, 8'd83, 8'd150, 8'd129, 8'd88, 8'd128, 8'd149, 8'd164, 8'd81, 8'd73, 8'd155, 8'd127, 8'd80, 8'd107, 8'd103, 8'd90, 8'd120, 8'd92, 8'd87, 8'd90, 8'd152, 8'd109, 8'd136, 8'd101, 8'd92, 8'd131, 8'd155, 8'd172, 8'd113, 8'd144, 8'd75, 8'd102, 8'd142, 8'd153, 8'd172, 8'd145, 8'd156, 8'd150, 8'd117, 8'd108, 8'd100, 8'd80, 8'd122, 8'd151, 8'd109, 8'd157, 8'd172, 8'd104, 8'd144, 8'd79, 8'd82, 8'd117, 8'd133, 8'd140, 8'd107, 8'd108, 8'd145, 8'd116, 8'd115, 8'd104, 8'd105, 8'd125, 8'd142, 8'd132, 8'd147, 8'd103, 8'd165, 8'd150, 8'd125, 8'd144, 8'd158, 8'd109, 8'd116, 8'd160, 8'd89, 8'd108, 8'd130, 8'd92, 8'd166, 8'd157, 8'd117, 8'd144, 8'd142, 8'd164, 8'd92, 8'd136, 8'd125, 8'd140, 8'd115, 8'd147, 8'd76, 8'd120, 8'd139, 8'd68, 8'd160, 8'd124, 8'd141, 8'd113, 8'd82, 8'd119, 8'd71, 8'd77, 8'd153, 8'd129, 8'd53, 8'd69, 8'd110, 8'd136, 8'd177, 8'd124, 8'd180, 8'd111, 8'd117, 8'd163, 8'd139, 8'd107, 8'd95, 8'd79, 8'd104, 8'd128, 8'd113, 8'd69, 8'd100, 8'd132, 8'd78, 8'd122, 8'd124, 8'd66, 8'd128, 8'd87, 8'd120, 8'd127, 8'd145, 8'd82, 8'd157, 8'd160, 8'd150, 8'd89, 8'd90, 8'd140, 8'd97, 8'd107, 8'd103, 8'd146, 8'd139, 8'd96, 8'd75, 8'd131, 8'd74, 8'd143, 8'd164, 8'd88, 8'd129, 8'd125, 8'd123, 8'd124, 8'd129, 8'd120, 8'd68, 8'd106, 8'd69, 8'd93, 8'd101, 8'd105, 8'd98, 8'd92, 8'd122, 8'd87, 8'd164, 8'd153, 8'd138, 8'd142, 8'd121, 8'd67, 8'd153, 8'd161, 8'd160, 8'd143, 8'd102, 8'd120, 8'd149, 8'd97, 8'd162, 8'd93, 8'd105, 8'd85, 8'd92, 8'd63, 8'd57, 8'd152, 8'd116, 8'd152, 8'd154, 8'd145, 8'd123, 8'd165, 8'd129, 8'd98, 8'd162, 8'd101, 8'd134, 8'd98, 8'd90, 8'd97, 8'd80, 8'd97, 8'd113, 8'd191, 8'd130, 8'd155, 8'd158, 8'd53, 8'd120, 8'd128, 8'd85, 8'd120, 8'd111, 8'd93, 8'd121, 8'd100, 8'd140, 8'd114, 8'd75, 8'd129, 8'd97, 8'd161, 8'd168, 8'd182, 8'd146, 8'd85, 8'd128, 8'd158, 8'd176, 8'd158, 8'd94, 8'd116, 8'd135, 8'd128, 8'd127, 8'd64, 8'd67, 8'd110, 8'd87, 8'd95, 8'd63, 8'd72, 8'd122, 8'd123, 8'd100, 8'd104, 8'd118, 8'd130, 8'd89, 8'd101, 8'd156, 8'd182, 8'd122, 8'd139, 8'd125, 8'd129, 8'd172, 8'd147, 8'd95, 8'd112, 8'd189, 8'd171, 8'd76, 8'd67, 8'd128, 8'd84, 8'd81, 8'd114, 8'd69, 8'd88, 8'd101, 8'd119, 8'd141, 8'd157, 8'd123, 8'd114, 8'd113, 8'd93, 8'd69, 8'd101, 8'd99, 8'd133, 8'd192, 8'd178, 8'd103, 8'd106, 8'd88, 8'd147, 8'd171, 8'd164, 8'd137, 8'd99, 8'd62, 8'd82, 8'd64, 8'd96, 8'd157, 8'd154, 8'd106, 8'd152, 8'd111, 8'd101, 8'd89, 8'd143, 8'd121, 8'd82, 8'd83, 8'd106, 8'd91, 8'd108, 8'd121, 8'd126, 8'd164, 8'd109, 8'd141, 8'd112, 8'd161, 8'd78, 8'd123, 8'd142, 8'd64, 8'd115, 8'd140, 8'd101, 8'd140, 8'd127, 8'd93, 8'd166, 8'd82, 8'd100, 8'd174, 8'd62, 8'd59, 8'd85, 8'd33, 8'd117, 8'd84, 8'd115, 8'd131, 8'd172, 8'd93, 8'd126, 8'd137, 8'd120, 8'd127, 8'd81, 8'd101, 8'd73, 8'd123, 8'd89, 8'd124, 8'd114, 8'd182, 8'd104, 8'd103, 8'd145, 8'd81, 8'd120, 8'd140, 8'd154, 8'd105, 8'd64, 8'd95, 8'd73, 8'd119, 8'd141, 8'd128, 8'd142, 8'd157, 8'd134, 8'd108, 8'd173, 8'd158, 8'd86, 8'd128, 8'd161, 8'd92, 8'd134, 8'd137, 8'd138, 8'd120, 8'd100, 8'd106, 8'd133, 8'd123, 8'd90, 8'd138, 8'd132, 8'd88, 8'd48, 8'd35, 8'd50, 8'd62, 8'd110, 8'd109, 8'd165, 8'd141, 8'd114, 8'd110, 8'd187, 8'd155, 8'd117, 8'd86, 8'd129, 8'd98, 8'd97, 8'd167, 8'd125, 8'd81, 8'd85, 8'd155, 8'd126, 8'd108, 8'd109, 8'd138, 8'd99, 8'd140, 8'd102, 8'd57, 8'd99, 8'd61, 8'd89, 8'd115, 8'd96, 8'd125, 8'd167, 8'd144, 8'd117, 8'd98, 8'd123, 8'd153, 8'd155, 8'd91, 8'd75, 8'd83, 8'd88, 8'd170, 8'd146, 8'd133, 8'd140, 8'd149, 8'd165, 8'd80, 8'd139, 8'd90, 8'd99, 8'd81, 8'd126, 8'd82, 8'd62, 8'd132, 8'd133, 8'd142, 8'd81, 8'd142, 8'd159, 8'd170, 8'd103, 8'd81, 8'd143, 8'd149, 8'd123, 8'd138, 8'd88, 8'd167, 8'd129, 8'd190, 8'd106, 8'd125, 8'd120, 8'd122, 8'd130, 8'd123, 8'd54, 8'd139, 8'd87, 8'd130, 8'd130, 8'd155, 8'd82, 8'd81, 8'd157, 8'd105, 8'd148, 8'd126, 8'd138, 8'd138, 8'd93, 8'd150, 8'd143, 8'd88, 8'd116, 8'd154, 8'd132, 8'd174, 8'd97, 8'd117, 8'd90, 8'd102, 8'd88, 8'd109, 8'd129, 8'd75, 8'd162, 8'd75, 8'd123, 8'd117, 8'd115, 8'd63, 8'd136, 8'd169, 8'd174, 8'd138, 8'd125, 8'd154, 8'd173, 8'd131, 8'd127, 8'd154, 8'd114, 8'd171, 8'd175, 8'd155, 8'd177, 8'd78, 8'd94, 8'd142, 8'd122, 8'd134, 8'd144, 8'd129, 8'd158, 8'd147, 8'd163, 8'd92, 8'd130, 8'd132, 8'd121, 8'd164, 8'd144, 8'd167, 8'd155, 8'd157, 8'd155, 8'd194, 8'd121, 8'd168, 8'd129, 8'd108, 8'd91, 8'd170, 8'd132, 8'd80, 8'd145, 8'd134, 8'd117, 8'd142, 8'd155, 8'd143, 8'd117, 8'd177, 8'd108, 8'd137, 8'd146, 8'd127, 8'd157, 8'd94, 8'd114, 8'd149, 8'd165, 8'd146, 8'd167, 8'd152, 8'd89, 8'd152, 8'd163, 8'd121, 8'd124, 8'd133, 8'd121, 8'd137, 8'd128, 8'd86, 8'd160, 8'd86, 8'd156, 8'd156, 8'd79, 8'd163, 8'd127, 8'd109, 8'd135, 8'd91, 8'd168, 8'd107, 8'd133, 8'd76, 8'd107, 8'd139, 8'd90, 8'd98, 8'd135, 8'd161, 8'd154, 8'd129, 8'd80, 8'd156, 8'd98, 8'd133, 8'd142, 8'd164})
) cell_0_6 (
    .clk(clk),
    .input_index(index_0_5_6),
    .input_value(value_0_5_6),
    .input_result(result_0_5_6),
    .input_enable(enable_0_5_6),
    .output_index(index_0_6_7),
    .output_value(value_0_6_7),
    .output_result(result_0_6_7),
    .output_enable(enable_0_6_7)
);

wire [10-1:0] index_0_7_8;
wire [`DATA_WIDTH-1:0] value_0_7_8;
wire [`DATA_WIDTH*4:0] result_0_7_8;
wire enable_0_7_8;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd114, 8'd141, 8'd99, 8'd114, 8'd110, 8'd108, 8'd84, 8'd137, 8'd113, 8'd87, 8'd61, 8'd99, 8'd93, 8'd81, 8'd119, 8'd148, 8'd157, 8'd130, 8'd92, 8'd147, 8'd129, 8'd133, 8'd133, 8'd121, 8'd73, 8'd167, 8'd123, 8'd96, 8'd101, 8'd166, 8'd122, 8'd156, 8'd109, 8'd155, 8'd136, 8'd145, 8'd101, 8'd125, 8'd60, 8'd60, 8'd31, 8'd46, 8'd133, 8'd129, 8'd97, 8'd50, 8'd110, 8'd55, 8'd63, 8'd132, 8'd148, 8'd81, 8'd87, 8'd101, 8'd109, 8'd139, 8'd70, 8'd106, 8'd122, 8'd134, 8'd140, 8'd130, 8'd60, 8'd88, 8'd86, 8'd147, 8'd72, 8'd80, 8'd102, 8'd140, 8'd87, 8'd107, 8'd80, 8'd137, 8'd93, 8'd112, 8'd88, 8'd95, 8'd63, 8'd90, 8'd119, 8'd125, 8'd149, 8'd118, 8'd109, 8'd146, 8'd152, 8'd159, 8'd96, 8'd76, 8'd104, 8'd64, 8'd135, 8'd141, 8'd105, 8'd80, 8'd169, 8'd119, 8'd152, 8'd151, 8'd137, 8'd105, 8'd94, 8'd145, 8'd61, 8'd86, 8'd94, 8'd159, 8'd142, 8'd166, 8'd116, 8'd93, 8'd79, 8'd165, 8'd125, 8'd170, 8'd145, 8'd154, 8'd167, 8'd165, 8'd101, 8'd96, 8'd137, 8'd116, 8'd94, 8'd105, 8'd92, 8'd150, 8'd145, 8'd145, 8'd123, 8'd135, 8'd139, 8'd137, 8'd92, 8'd180, 8'd179, 8'd134, 8'd124, 8'd95, 8'd158, 8'd131, 8'd129, 8'd92, 8'd132, 8'd177, 8'd129, 8'd151, 8'd130, 8'd139, 8'd134, 8'd88, 8'd173, 8'd116, 8'd185, 8'd163, 8'd186, 8'd134, 8'd123, 8'd119, 8'd157, 8'd122, 8'd93, 8'd133, 8'd112, 8'd123, 8'd134, 8'd92, 8'd156, 8'd133, 8'd123, 8'd154, 8'd117, 8'd112, 8'd190, 8'd153, 8'd135, 8'd103, 8'd99, 8'd150, 8'd107, 8'd140, 8'd172, 8'd147, 8'd138, 8'd112, 8'd144, 8'd154, 8'd140, 8'd137, 8'd101, 8'd131, 8'd116, 8'd112, 8'd164, 8'd87, 8'd103, 8'd106, 8'd161, 8'd172, 8'd125, 8'd176, 8'd132, 8'd153, 8'd179, 8'd155, 8'd114, 8'd127, 8'd184, 8'd152, 8'd112, 8'd121, 8'd107, 8'd144, 8'd113, 8'd186, 8'd121, 8'd124, 8'd162, 8'd121, 8'd191, 8'd164, 8'd157, 8'd129, 8'd76, 8'd172, 8'd133, 8'd145, 8'd172, 8'd194, 8'd195, 8'd141, 8'd184, 8'd193, 8'd118, 8'd140, 8'd94, 8'd82, 8'd89, 8'd150, 8'd163, 8'd119, 8'd148, 8'd132, 8'd118, 8'd138, 8'd153, 8'd141, 8'd171, 8'd172, 8'd140, 8'd127, 8'd169, 8'd103, 8'd108, 8'd200, 8'd147, 8'd189, 8'd137, 8'd189, 8'd119, 8'd171, 8'd110, 8'd144, 8'd149, 8'd122, 8'd114, 8'd169, 8'd173, 8'd105, 8'd99, 8'd167, 8'd117, 8'd166, 8'd144, 8'd178, 8'd145, 8'd86, 8'd125, 8'd114, 8'd174, 8'd134, 8'd178, 8'd111, 8'd195, 8'd166, 8'd187, 8'd166, 8'd90, 8'd91, 8'd85, 8'd167, 8'd121, 8'd134, 8'd59, 8'd163, 8'd134, 8'd118, 8'd159, 8'd132, 8'd74, 8'd164, 8'd116, 8'd146, 8'd189, 8'd84, 8'd134, 8'd95, 8'd141, 8'd118, 8'd191, 8'd134, 8'd143, 8'd123, 8'd159, 8'd95, 8'd158, 8'd113, 8'd59, 8'd113, 8'd91, 8'd153, 8'd79, 8'd100, 8'd176, 8'd105, 8'd136, 8'd147, 8'd87, 8'd67, 8'd111, 8'd108, 8'd166, 8'd142, 8'd151, 8'd77, 8'd119, 8'd163, 8'd114, 8'd122, 8'd93, 8'd103, 8'd101, 8'd135, 8'd91, 8'd105, 8'd123, 8'd129, 8'd125, 8'd109, 8'd164, 8'd179, 8'd148, 8'd198, 8'd113, 8'd118, 8'd145, 8'd146, 8'd80, 8'd108, 8'd134, 8'd149, 8'd83, 8'd94, 8'd123, 8'd176, 8'd172, 8'd116, 8'd140, 8'd156, 8'd128, 8'd66, 8'd100, 8'd85, 8'd123, 8'd111, 8'd98, 8'd97, 8'd104, 8'd171, 8'd187, 8'd155, 8'd159, 8'd141, 8'd116, 8'd76, 8'd51, 8'd95, 8'd128, 8'd56, 8'd100, 8'd168, 8'd86, 8'd173, 8'd118, 8'd123, 8'd147, 8'd124, 8'd52, 8'd102, 8'd123, 8'd138, 8'd88, 8'd65, 8'd123, 8'd110, 8'd127, 8'd143, 8'd155, 8'd152, 8'd89, 8'd131, 8'd83, 8'd76, 8'd143, 8'd74, 8'd139, 8'd107, 8'd156, 8'd156, 8'd139, 8'd169, 8'd186, 8'd94, 8'd53, 8'd123, 8'd30, 8'd69, 8'd113, 8'd55, 8'd55, 8'd133, 8'd90, 8'd139, 8'd126, 8'd154, 8'd157, 8'd86, 8'd100, 8'd108, 8'd91, 8'd98, 8'd125, 8'd116, 8'd93, 8'd77, 8'd108, 8'd123, 8'd144, 8'd157, 8'd193, 8'd197, 8'd119, 8'd100, 8'd37, 8'd77, 8'd85, 8'd123, 8'd116, 8'd112, 8'd30, 8'd65, 8'd121, 8'd153, 8'd111, 8'd122, 8'd111, 8'd108, 8'd146, 8'd116, 8'd106, 8'd99, 8'd105, 8'd139, 8'd75, 8'd142, 8'd138, 8'd191, 8'd168, 8'd190, 8'd206, 8'd128, 8'd71, 8'd126, 8'd65, 8'd51, 8'd98, 8'd118, 8'd76, 8'd121, 8'd116, 8'd113, 8'd148, 8'd129, 8'd146, 8'd139, 8'd153, 8'd91, 8'd66, 8'd118, 8'd72, 8'd63, 8'd134, 8'd114, 8'd128, 8'd142, 8'd136, 8'd199, 8'd153, 8'd133, 8'd82, 8'd107, 8'd126, 8'd77, 8'd41, 8'd113, 8'd96, 8'd128, 8'd153, 8'd128, 8'd142, 8'd140, 8'd72, 8'd129, 8'd124, 8'd118, 8'd62, 8'd74, 8'd72, 8'd120, 8'd71, 8'd132, 8'd146, 8'd164, 8'd203, 8'd158, 8'd142, 8'd172, 8'd171, 8'd86, 8'd121, 8'd122, 8'd130, 8'd124, 8'd67, 8'd115, 8'd72, 8'd108, 8'd156, 8'd155, 8'd114, 8'd131, 8'd65, 8'd82, 8'd149, 8'd147, 8'd117, 8'd147, 8'd120, 8'd81, 8'd175, 8'd88, 8'd214, 8'd175, 8'd104, 8'd166, 8'd166, 8'd156, 8'd84, 8'd99, 8'd95, 8'd129, 8'd79, 8'd135, 8'd163, 8'd141, 8'd91, 8'd73, 8'd83, 8'd77, 8'd122, 8'd74, 8'd112, 8'd155, 8'd96, 8'd138, 8'd103, 8'd120, 8'd153, 8'd189, 8'd153, 8'd139, 8'd149, 8'd165, 8'd168, 8'd144, 8'd106, 8'd144, 8'd138, 8'd174, 8'd171, 8'd162, 8'd90, 8'd142, 8'd122, 8'd145, 8'd92, 8'd114, 8'd88, 8'd111, 8'd116, 8'd91, 8'd139, 8'd117, 8'd90, 8'd154, 8'd160, 8'd126, 8'd147, 8'd158, 8'd114, 8'd158, 8'd150, 8'd111, 8'd163, 8'd154, 8'd169, 8'd178, 8'd98, 8'd141, 8'd91, 8'd94, 8'd142, 8'd141, 8'd170, 8'd157, 8'd138, 8'd128, 8'd126, 8'd158, 8'd125, 8'd158, 8'd154, 8'd97, 8'd91, 8'd159, 8'd174, 8'd156, 8'd165, 8'd82, 8'd99, 8'd98, 8'd93, 8'd111, 8'd116, 8'd164, 8'd113, 8'd173, 8'd135, 8'd162, 8'd119, 8'd122, 8'd166, 8'd171, 8'd180, 8'd99, 8'd132, 8'd145, 8'd129, 8'd153, 8'd164, 8'd96, 8'd77, 8'd113, 8'd116, 8'd103, 8'd78, 8'd100, 8'd167, 8'd136, 8'd110, 8'd151, 8'd130, 8'd140, 8'd124, 8'd207, 8'd136, 8'd136, 8'd210, 8'd203, 8'd173, 8'd121, 8'd94, 8'd98, 8'd167, 8'd149, 8'd107, 8'd153, 8'd124, 8'd84, 8'd84, 8'd148, 8'd114, 8'd130, 8'd78, 8'd79, 8'd71, 8'd91, 8'd186, 8'd152, 8'd142, 8'd112, 8'd106, 8'd152, 8'd126, 8'd127, 8'd166, 8'd188, 8'd127, 8'd156, 8'd108, 8'd153, 8'd106, 8'd76, 8'd148, 8'd94, 8'd109, 8'd153, 8'd115, 8'd134, 8'd148, 8'd148, 8'd119, 8'd129, 8'd81, 8'd132, 8'd183, 8'd172, 8'd144, 8'd185, 8'd78, 8'd150, 8'd155, 8'd103, 8'd152, 8'd103, 8'd122, 8'd136, 8'd108, 8'd141, 8'd165, 8'd138, 8'd159, 8'd74, 8'd113, 8'd143, 8'd119, 8'd120, 8'd144, 8'd168, 8'd103, 8'd155, 8'd135, 8'd78, 8'd71, 8'd127, 8'd136, 8'd77, 8'd105, 8'd74, 8'd78, 8'd175, 8'd97, 8'd142, 8'd142, 8'd111, 8'd88, 8'd126, 8'd94, 8'd103, 8'd155, 8'd136, 8'd120, 8'd165})
) cell_0_7 (
    .clk(clk),
    .input_index(index_0_6_7),
    .input_value(value_0_6_7),
    .input_result(result_0_6_7),
    .input_enable(enable_0_6_7),
    .output_index(index_0_7_8),
    .output_value(value_0_7_8),
    .output_result(result_0_7_8),
    .output_enable(enable_0_7_8)
);

wire [10-1:0] index_0_8_9;
wire [`DATA_WIDTH-1:0] value_0_8_9;
wire [`DATA_WIDTH*4:0] result_0_8_9;
wire enable_0_8_9;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd70, 8'd109, 8'd112, 8'd114, 8'd107, 8'd143, 8'd89, 8'd153, 8'd112, 8'd178, 8'd141, 8'd180, 8'd97, 8'd133, 8'd100, 8'd157, 8'd139, 8'd153, 8'd87, 8'd83, 8'd70, 8'd90, 8'd139, 8'd143, 8'd114, 8'd78, 8'd157, 8'd152, 8'd97, 8'd119, 8'd106, 8'd125, 8'd130, 8'd142, 8'd137, 8'd142, 8'd118, 8'd152, 8'd126, 8'd143, 8'd78, 8'd77, 8'd104, 8'd80, 8'd135, 8'd133, 8'd75, 8'd128, 8'd123, 8'd109, 8'd122, 8'd67, 8'd87, 8'd138, 8'd99, 8'd98, 8'd125, 8'd119, 8'd145, 8'd83, 8'd88, 8'd149, 8'd118, 8'd96, 8'd119, 8'd152, 8'd83, 8'd96, 8'd91, 8'd147, 8'd129, 8'd99, 8'd126, 8'd114, 8'd157, 8'd152, 8'd147, 8'd169, 8'd95, 8'd127, 8'd172, 8'd110, 8'd137, 8'd144, 8'd109, 8'd147, 8'd85, 8'd94, 8'd116, 8'd125, 8'd126, 8'd70, 8'd77, 8'd67, 8'd93, 8'd164, 8'd84, 8'd149, 8'd120, 8'd129, 8'd131, 8'd148, 8'd132, 8'd141, 8'd90, 8'd157, 8'd114, 8'd185, 8'd136, 8'd168, 8'd121, 8'd121, 8'd83, 8'd115, 8'd130, 8'd161, 8'd116, 8'd148, 8'd100, 8'd114, 8'd144, 8'd157, 8'd81, 8'd100, 8'd106, 8'd77, 8'd61, 8'd114, 8'd158, 8'd158, 8'd115, 8'd119, 8'd162, 8'd115, 8'd142, 8'd120, 8'd196, 8'd168, 8'd161, 8'd111, 8'd83, 8'd101, 8'd170, 8'd164, 8'd105, 8'd150, 8'd95, 8'd168, 8'd79, 8'd151, 8'd78, 8'd121, 8'd139, 8'd163, 8'd103, 8'd129, 8'd176, 8'd164, 8'd87, 8'd160, 8'd158, 8'd164, 8'd162, 8'd172, 8'd192, 8'd180, 8'd129, 8'd115, 8'd105, 8'd127, 8'd133, 8'd101, 8'd153, 8'd103, 8'd172, 8'd144, 8'd94, 8'd129, 8'd173, 8'd99, 8'd181, 8'd94, 8'd144, 8'd92, 8'd92, 8'd93, 8'd117, 8'd95, 8'd159, 8'd163, 8'd108, 8'd120, 8'd137, 8'd114, 8'd124, 8'd110, 8'd168, 8'd101, 8'd128, 8'd131, 8'd123, 8'd151, 8'd158, 8'd169, 8'd156, 8'd125, 8'd170, 8'd115, 8'd110, 8'd128, 8'd152, 8'd181, 8'd154, 8'd191, 8'd165, 8'd173, 8'd139, 8'd166, 8'd113, 8'd107, 8'd202, 8'd120, 8'd108, 8'd139, 8'd157, 8'd112, 8'd115, 8'd145, 8'd99, 8'd176, 8'd127, 8'd184, 8'd111, 8'd91, 8'd138, 8'd139, 8'd168, 8'd95, 8'd113, 8'd146, 8'd195, 8'd126, 8'd91, 8'd87, 8'd99, 8'd112, 8'd112, 8'd162, 8'd137, 8'd143, 8'd166, 8'd160, 8'd100, 8'd148, 8'd201, 8'd164, 8'd162, 8'd107, 8'd148, 8'd187, 8'd99, 8'd90, 8'd99, 8'd90, 8'd138, 8'd88, 8'd117, 8'd104, 8'd108, 8'd113, 8'd105, 8'd116, 8'd96, 8'd143, 8'd127, 8'd162, 8'd185, 8'd167, 8'd90, 8'd83, 8'd118, 8'd148, 8'd171, 8'd126, 8'd139, 8'd183, 8'd108, 8'd101, 8'd179, 8'd140, 8'd117, 8'd123, 8'd125, 8'd71, 8'd103, 8'd53, 8'd127, 8'd156, 8'd76, 8'd133, 8'd149, 8'd109, 8'd106, 8'd112, 8'd139, 8'd148, 8'd111, 8'd76, 8'd96, 8'd173, 8'd116, 8'd207, 8'd114, 8'd164, 8'd109, 8'd97, 8'd173, 8'd94, 8'd69, 8'd85, 8'd126, 8'd98, 8'd97, 8'd154, 8'd160, 8'd136, 8'd131, 8'd146, 8'd146, 8'd98, 8'd107, 8'd119, 8'd145, 8'd117, 8'd127, 8'd89, 8'd121, 8'd126, 8'd137, 8'd202, 8'd181, 8'd107, 8'd139, 8'd154, 8'd114, 8'd67, 8'd141, 8'd129, 8'd75, 8'd88, 8'd65, 8'd131, 8'd78, 8'd111, 8'd158, 8'd123, 8'd120, 8'd166, 8'd121, 8'd71, 8'd122, 8'd132, 8'd91, 8'd88, 8'd123, 8'd174, 8'd100, 8'd154, 8'd123, 8'd108, 8'd166, 8'd90, 8'd114, 8'd112, 8'd78, 8'd104, 8'd140, 8'd97, 8'd156, 8'd80, 8'd152, 8'd169, 8'd134, 8'd168, 8'd169, 8'd121, 8'd98, 8'd61, 8'd82, 8'd124, 8'd83, 8'd142, 8'd109, 8'd192, 8'd103, 8'd103, 8'd71, 8'd145, 8'd81, 8'd70, 8'd130, 8'd56, 8'd100, 8'd46, 8'd75, 8'd134, 8'd133, 8'd151, 8'd104, 8'd149, 8'd135, 8'd142, 8'd140, 8'd67, 8'd115, 8'd150, 8'd152, 8'd140, 8'd136, 8'd76, 8'd89, 8'd159, 8'd144, 8'd80, 8'd123, 8'd22, 8'd118, 8'd47, 8'd122, 8'd130, 8'd117, 8'd78, 8'd121, 8'd78, 8'd118, 8'd164, 8'd121, 8'd68, 8'd141, 8'd146, 8'd82, 8'd144, 8'd142, 8'd92, 8'd148, 8'd129, 8'd155, 8'd162, 8'd76, 8'd88, 8'd162, 8'd131, 8'd126, 8'd100, 8'd89, 8'd117, 8'd80, 8'd86, 8'd139, 8'd107, 8'd79, 8'd140, 8'd83, 8'd149, 8'd118, 8'd65, 8'd145, 8'd43, 8'd117, 8'd88, 8'd69, 8'd148, 8'd111, 8'd167, 8'd190, 8'd163, 8'd77, 8'd172, 8'd160, 8'd138, 8'd134, 8'd96, 8'd146, 8'd66, 8'd117, 8'd130, 8'd114, 8'd132, 8'd143, 8'd138, 8'd148, 8'd143, 8'd78, 8'd129, 8'd112, 8'd153, 8'd118, 8'd105, 8'd91, 8'd147, 8'd178, 8'd164, 8'd167, 8'd103, 8'd125, 8'd119, 8'd119, 8'd116, 8'd103, 8'd153, 8'd130, 8'd133, 8'd70, 8'd55, 8'd156, 8'd92, 8'd106, 8'd102, 8'd130, 8'd74, 8'd166, 8'd127, 8'd88, 8'd91, 8'd80, 8'd97, 8'd75, 8'd161, 8'd175, 8'd106, 8'd144, 8'd118, 8'd133, 8'd131, 8'd120, 8'd98, 8'd91, 8'd101, 8'd100, 8'd100, 8'd100, 8'd86, 8'd148, 8'd153, 8'd162, 8'd102, 8'd164, 8'd125, 8'd101, 8'd153, 8'd120, 8'd154, 8'd143, 8'd127, 8'd111, 8'd120, 8'd87, 8'd116, 8'd172, 8'd95, 8'd125, 8'd118, 8'd101, 8'd136, 8'd109, 8'd139, 8'd111, 8'd103, 8'd114, 8'd129, 8'd154, 8'd109, 8'd107, 8'd93, 8'd95, 8'd162, 8'd137, 8'd123, 8'd119, 8'd144, 8'd114, 8'd119, 8'd153, 8'd94, 8'd137, 8'd121, 8'd168, 8'd86, 8'd120, 8'd179, 8'd129, 8'd120, 8'd102, 8'd111, 8'd135, 8'd159, 8'd117, 8'd106, 8'd80, 8'd77, 8'd89, 8'd125, 8'd107, 8'd139, 8'd152, 8'd101, 8'd95, 8'd177, 8'd89, 8'd91, 8'd89, 8'd108, 8'd78, 8'd90, 8'd166, 8'd168, 8'd111, 8'd127, 8'd152, 8'd145, 8'd166, 8'd139, 8'd143, 8'd152, 8'd98, 8'd139, 8'd163, 8'd89, 8'd136, 8'd151, 8'd144, 8'd129, 8'd145, 8'd169, 8'd108, 8'd176, 8'd126, 8'd92, 8'd93, 8'd87, 8'd122, 8'd110, 8'd76, 8'd149, 8'd124, 8'd123, 8'd162, 8'd173, 8'd120, 8'd96, 8'd132, 8'd89, 8'd120, 8'd158, 8'd193, 8'd163, 8'd173, 8'd146, 8'd158, 8'd162, 8'd122, 8'd152, 8'd153, 8'd168, 8'd109, 8'd169, 8'd149, 8'd160, 8'd145, 8'd98, 8'd154, 8'd130, 8'd88, 8'd84, 8'd117, 8'd168, 8'd150, 8'd102, 8'd177, 8'd141, 8'd160, 8'd147, 8'd131, 8'd203, 8'd129, 8'd203, 8'd156, 8'd157, 8'd228, 8'd170, 8'd166, 8'd195, 8'd197, 8'd180, 8'd159, 8'd164, 8'd158, 8'd70, 8'd72, 8'd161, 8'd113, 8'd112, 8'd163, 8'd92, 8'd157, 8'd132, 8'd162, 8'd134, 8'd155, 8'd136, 8'd175, 8'd140, 8'd162, 8'd127, 8'd111, 8'd154, 8'd211, 8'd199, 8'd144, 8'd185, 8'd135, 8'd141, 8'd76, 8'd92, 8'd106, 8'd139, 8'd169, 8'd119, 8'd102, 8'd81, 8'd145, 8'd113, 8'd152, 8'd171, 8'd151, 8'd124, 8'd185, 8'd102, 8'd161, 8'd133, 8'd151, 8'd138, 8'd199, 8'd185, 8'd189, 8'd181, 8'd172, 8'd125, 8'd133, 8'd147, 8'd98, 8'd161, 8'd110, 8'd90, 8'd95, 8'd72, 8'd159, 8'd100, 8'd154, 8'd122, 8'd77, 8'd76, 8'd93, 8'd71, 8'd138, 8'd103, 8'd104, 8'd101, 8'd102, 8'd92, 8'd155, 8'd142, 8'd163, 8'd98, 8'd98, 8'd83, 8'd169, 8'd124, 8'd164, 8'd137, 8'd140, 8'd120, 8'd152, 8'd153})
) cell_0_8 (
    .clk(clk),
    .input_index(index_0_7_8),
    .input_value(value_0_7_8),
    .input_result(result_0_7_8),
    .input_enable(enable_0_7_8),
    .output_index(index_0_8_9),
    .output_value(value_0_8_9),
    .output_result(result_0_8_9),
    .output_enable(enable_0_8_9)
);

wire [10-1:0] index_0_9_10;
wire [`DATA_WIDTH-1:0] value_0_9_10;
wire [`DATA_WIDTH*4:0] result_0_9_10;
wire enable_0_9_10;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd77, 8'd124, 8'd164, 8'd129, 8'd148, 8'd78, 8'd100, 8'd143, 8'd112, 8'd133, 8'd61, 8'd80, 8'd85, 8'd104, 8'd65, 8'd111, 8'd93, 8'd114, 8'd78, 8'd85, 8'd102, 8'd88, 8'd133, 8'd129, 8'd139, 8'd128, 8'd161, 8'd164, 8'd162, 8'd111, 8'd80, 8'd78, 8'd142, 8'd76, 8'd68, 8'd77, 8'd38, 8'd121, 8'd118, 8'd71, 8'd81, 8'd23, 8'd68, 8'd25, 8'd65, 8'd51, 8'd49, 8'd107, 8'd57, 8'd52, 8'd76, 8'd142, 8'd82, 8'd100, 8'd72, 8'd150, 8'd160, 8'd111, 8'd166, 8'd155, 8'd109, 8'd157, 8'd124, 8'd105, 8'd66, 8'd128, 8'd122, 8'd97, 8'd143, 8'd101, 8'd129, 8'd96, 8'd43, 8'd84, 8'd90, 8'd120, 8'd135, 8'd138, 8'd107, 8'd116, 8'd161, 8'd168, 8'd72, 8'd95, 8'd80, 8'd144, 8'd129, 8'd88, 8'd115, 8'd142, 8'd71, 8'd84, 8'd67, 8'd138, 8'd154, 8'd126, 8'd64, 8'd74, 8'd151, 8'd101, 8'd85, 8'd77, 8'd140, 8'd104, 8'd62, 8'd59, 8'd69, 8'd117, 8'd125, 8'd109, 8'd101, 8'd106, 8'd72, 8'd101, 8'd134, 8'd114, 8'd101, 8'd136, 8'd132, 8'd96, 8'd101, 8'd95, 8'd68, 8'd137, 8'd137, 8'd69, 8'd116, 8'd92, 8'd117, 8'd80, 8'd113, 8'd84, 8'd93, 8'd113, 8'd146, 8'd173, 8'd188, 8'd133, 8'd149, 8'd133, 8'd145, 8'd82, 8'd145, 8'd165, 8'd89, 8'd105, 8'd158, 8'd163, 8'd164, 8'd152, 8'd94, 8'd93, 8'd119, 8'd132, 8'd138, 8'd109, 8'd136, 8'd169, 8'd106, 8'd118, 8'd72, 8'd68, 8'd160, 8'd161, 8'd124, 8'd130, 8'd102, 8'd81, 8'd169, 8'd178, 8'd91, 8'd135, 8'd173, 8'd183, 8'd166, 8'd161, 8'd116, 8'd103, 8'd126, 8'd85, 8'd125, 8'd92, 8'd89, 8'd107, 8'd139, 8'd92, 8'd138, 8'd102, 8'd91, 8'd86, 8'd159, 8'd135, 8'd166, 8'd159, 8'd99, 8'd65, 8'd72, 8'd158, 8'd137, 8'd101, 8'd177, 8'd130, 8'd108, 8'd151, 8'd137, 8'd94, 8'd114, 8'd158, 8'd105, 8'd180, 8'd107, 8'd123, 8'd130, 8'd194, 8'd109, 8'd161, 8'd84, 8'd146, 8'd97, 8'd119, 8'd127, 8'd138, 8'd139, 8'd106, 8'd150, 8'd129, 8'd175, 8'd102, 8'd166, 8'd87, 8'd168, 8'd144, 8'd128, 8'd155, 8'd86, 8'd130, 8'd98, 8'd102, 8'd140, 8'd127, 8'd109, 8'd151, 8'd109, 8'd171, 8'd173, 8'd99, 8'd139, 8'd128, 8'd91, 8'd85, 8'd141, 8'd70, 8'd142, 8'd88, 8'd155, 8'd192, 8'd134, 8'd162, 8'd161, 8'd89, 8'd124, 8'd130, 8'd125, 8'd107, 8'd148, 8'd172, 8'd116, 8'd138, 8'd111, 8'd117, 8'd108, 8'd140, 8'd164, 8'd119, 8'd174, 8'd150, 8'd131, 8'd95, 8'd152, 8'd130, 8'd117, 8'd104, 8'd200, 8'd105, 8'd183, 8'd155, 8'd150, 8'd159, 8'd115, 8'd145, 8'd163, 8'd155, 8'd75, 8'd152, 8'd161, 8'd85, 8'd123, 8'd135, 8'd96, 8'd150, 8'd114, 8'd187, 8'd119, 8'd129, 8'd146, 8'd108, 8'd147, 8'd164, 8'd128, 8'd186, 8'd173, 8'd183, 8'd103, 8'd175, 8'd156, 8'd110, 8'd97, 8'd153, 8'd130, 8'd150, 8'd84, 8'd116, 8'd157, 8'd109, 8'd144, 8'd157, 8'd94, 8'd159, 8'd104, 8'd123, 8'd127, 8'd90, 8'd66, 8'd114, 8'd149, 8'd88, 8'd158, 8'd204, 8'd175, 8'd163, 8'd172, 8'd150, 8'd87, 8'd88, 8'd84, 8'd140, 8'd63, 8'd115, 8'd81, 8'd83, 8'd103, 8'd142, 8'd201, 8'd195, 8'd197, 8'd148, 8'd109, 8'd131, 8'd100, 8'd107, 8'd61, 8'd117, 8'd147, 8'd89, 8'd138, 8'd141, 8'd183, 8'd161, 8'd152, 8'd159, 8'd130, 8'd111, 8'd140, 8'd66, 8'd106, 8'd82, 8'd130, 8'd88, 8'd115, 8'd170, 8'd137, 8'd157, 8'd169, 8'd137, 8'd184, 8'd124, 8'd102, 8'd138, 8'd106, 8'd152, 8'd149, 8'd158, 8'd125, 8'd114, 8'd105, 8'd161, 8'd143, 8'd86, 8'd161, 8'd122, 8'd78, 8'd66, 8'd66, 8'd86, 8'd73, 8'd63, 8'd109, 8'd185, 8'd163, 8'd123, 8'd133, 8'd100, 8'd144, 8'd147, 8'd132, 8'd51, 8'd100, 8'd79, 8'd114, 8'd76, 8'd167, 8'd172, 8'd177, 8'd149, 8'd142, 8'd140, 8'd97, 8'd94, 8'd128, 8'd99, 8'd95, 8'd138, 8'd42, 8'd90, 8'd78, 8'd99, 8'd164, 8'd167, 8'd136, 8'd91, 8'd87, 8'd65, 8'd116, 8'd96, 8'd60, 8'd121, 8'd141, 8'd156, 8'd167, 8'd105, 8'd126, 8'd167, 8'd118, 8'd77, 8'd71, 8'd117, 8'd107, 8'd70, 8'd80, 8'd51, 8'd63, 8'd61, 8'd106, 8'd161, 8'd110, 8'd123, 8'd74, 8'd107, 8'd79, 8'd55, 8'd58, 8'd61, 8'd129, 8'd55, 8'd85, 8'd135, 8'd147, 8'd102, 8'd128, 8'd210, 8'd149, 8'd137, 8'd85, 8'd133, 8'd148, 8'd110, 8'd69, 8'd122, 8'd48, 8'd47, 8'd150, 8'd108, 8'd97, 8'd136, 8'd82, 8'd141, 8'd103, 8'd146, 8'd140, 8'd137, 8'd81, 8'd132, 8'd140, 8'd85, 8'd122, 8'd167, 8'd150, 8'd195, 8'd154, 8'd165, 8'd120, 8'd147, 8'd134, 8'd78, 8'd78, 8'd138, 8'd75, 8'd80, 8'd119, 8'd141, 8'd144, 8'd114, 8'd107, 8'd145, 8'd117, 8'd127, 8'd157, 8'd108, 8'd117, 8'd69, 8'd127, 8'd128, 8'd145, 8'd106, 8'd134, 8'd137, 8'd98, 8'd99, 8'd75, 8'd74, 8'd135, 8'd71, 8'd142, 8'd119, 8'd79, 8'd114, 8'd137, 8'd113, 8'd150, 8'd123, 8'd165, 8'd89, 8'd146, 8'd65, 8'd141, 8'd133, 8'd141, 8'd90, 8'd147, 8'd113, 8'd118, 8'd164, 8'd152, 8'd156, 8'd109, 8'd180, 8'd139, 8'd142, 8'd63, 8'd126, 8'd125, 8'd145, 8'd62, 8'd87, 8'd71, 8'd71, 8'd123, 8'd98, 8'd126, 8'd104, 8'd119, 8'd159, 8'd90, 8'd140, 8'd80, 8'd97, 8'd118, 8'd145, 8'd90, 8'd104, 8'd146, 8'd124, 8'd103, 8'd131, 8'd119, 8'd111, 8'd139, 8'd164, 8'd83, 8'd120, 8'd140, 8'd99, 8'd59, 8'd126, 8'd147, 8'd126, 8'd169, 8'd80, 8'd125, 8'd76, 8'd107, 8'd176, 8'd84, 8'd153, 8'd123, 8'd132, 8'd176, 8'd180, 8'd93, 8'd183, 8'd102, 8'd105, 8'd110, 8'd109, 8'd182, 8'd179, 8'd201, 8'd110, 8'd126, 8'd95, 8'd94, 8'd158, 8'd85, 8'd179, 8'd151, 8'd169, 8'd138, 8'd121, 8'd135, 8'd149, 8'd108, 8'd126, 8'd119, 8'd104, 8'd155, 8'd138, 8'd101, 8'd131, 8'd133, 8'd137, 8'd100, 8'd131, 8'd173, 8'd131, 8'd151, 8'd147, 8'd108, 8'd88, 8'd165, 8'd182, 8'd182, 8'd87, 8'd178, 8'd142, 8'd104, 8'd105, 8'd117, 8'd121, 8'd119, 8'd86, 8'd113, 8'd145, 8'd81, 8'd137, 8'd97, 8'd128, 8'd141, 8'd161, 8'd114, 8'd195, 8'd164, 8'd193, 8'd142, 8'd143, 8'd128, 8'd132, 8'd165, 8'd113, 8'd159, 8'd171, 8'd113, 8'd130, 8'd90, 8'd133, 8'd150, 8'd103, 8'd116, 8'd130, 8'd98, 8'd139, 8'd127, 8'd166, 8'd151, 8'd167, 8'd130, 8'd107, 8'd128, 8'd168, 8'd179, 8'd177, 8'd120, 8'd167, 8'd157, 8'd100, 8'd72, 8'd124, 8'd92, 8'd174, 8'd162, 8'd149, 8'd69, 8'd103, 8'd157, 8'd95, 8'd96, 8'd74, 8'd145, 8'd151, 8'd148, 8'd87, 8'd161, 8'd142, 8'd128, 8'd118, 8'd78, 8'd90, 8'd87, 8'd154, 8'd171, 8'd109, 8'd122, 8'd144, 8'd145, 8'd115, 8'd100, 8'd86, 8'd112, 8'd112, 8'd80, 8'd62, 8'd129, 8'd77, 8'd123, 8'd124, 8'd82, 8'd123, 8'd80, 8'd107, 8'd170, 8'd101, 8'd83, 8'd132, 8'd85, 8'd155, 8'd71, 8'd81, 8'd89, 8'd121, 8'd147, 8'd90, 8'd81, 8'd161, 8'd169, 8'd89, 8'd137, 8'd90, 8'd101, 8'd132, 8'd127, 8'd168, 8'd168, 8'd123, 8'd105, 8'd165})
) cell_0_9 (
    .clk(clk),
    .input_index(index_0_8_9),
    .input_value(value_0_8_9),
    .input_result(result_0_8_9),
    .input_enable(enable_0_8_9),
    .output_index(index_0_9_10),
    .output_value(value_0_9_10),
    .output_result(result_0_9_10),
    .output_enable(enable_0_9_10)
);

wire [10-1:0] index_0_10_11;
wire [`DATA_WIDTH-1:0] value_0_10_11;
wire [`DATA_WIDTH*4:0] result_0_10_11;
wire enable_0_10_11;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd153, 8'd151, 8'd102, 8'd84, 8'd100, 8'd128, 8'd179, 8'd113, 8'd177, 8'd100, 8'd90, 8'd162, 8'd194, 8'd191, 8'd169, 8'd94, 8'd77, 8'd89, 8'd157, 8'd179, 8'd168, 8'd118, 8'd125, 8'd112, 8'd149, 8'd122, 8'd136, 8'd130, 8'd114, 8'd106, 8'd147, 8'd109, 8'd130, 8'd121, 8'd157, 8'd155, 8'd162, 8'd143, 8'd147, 8'd155, 8'd188, 8'd160, 8'd104, 8'd153, 8'd156, 8'd101, 8'd186, 8'd153, 8'd194, 8'd123, 8'd144, 8'd154, 8'd138, 8'd152, 8'd110, 8'd116, 8'd109, 8'd105, 8'd158, 8'd126, 8'd108, 8'd123, 8'd110, 8'd175, 8'd88, 8'd155, 8'd123, 8'd140, 8'd157, 8'd82, 8'd143, 8'd159, 8'd113, 8'd150, 8'd137, 8'd153, 8'd148, 8'd116, 8'd95, 8'd115, 8'd106, 8'd91, 8'd158, 8'd81, 8'd75, 8'd154, 8'd130, 8'd152, 8'd116, 8'd107, 8'd134, 8'd165, 8'd169, 8'd109, 8'd129, 8'd107, 8'd155, 8'd105, 8'd124, 8'd74, 8'd128, 8'd150, 8'd103, 8'd155, 8'd158, 8'd140, 8'd143, 8'd138, 8'd135, 8'd146, 8'd126, 8'd77, 8'd147, 8'd110, 8'd96, 8'd97, 8'd115, 8'd76, 8'd160, 8'd121, 8'd114, 8'd111, 8'd151, 8'd109, 8'd111, 8'd167, 8'd124, 8'd130, 8'd93, 8'd94, 8'd139, 8'd165, 8'd128, 8'd109, 8'd142, 8'd144, 8'd103, 8'd56, 8'd158, 8'd104, 8'd93, 8'd150, 8'd125, 8'd163, 8'd134, 8'd66, 8'd115, 8'd100, 8'd121, 8'd98, 8'd163, 8'd108, 8'd91, 8'd133, 8'd96, 8'd103, 8'd93, 8'd111, 8'd91, 8'd118, 8'd131, 8'd163, 8'd77, 8'd81, 8'd118, 8'd151, 8'd163, 8'd158, 8'd130, 8'd61, 8'd94, 8'd150, 8'd113, 8'd87, 8'd63, 8'd92, 8'd144, 8'd98, 8'd112, 8'd147, 8'd157, 8'd121, 8'd132, 8'd78, 8'd142, 8'd93, 8'd130, 8'd100, 8'd96, 8'd103, 8'd112, 8'd56, 8'd113, 8'd72, 8'd97, 8'd119, 8'd82, 8'd162, 8'd118, 8'd113, 8'd91, 8'd73, 8'd81, 8'd78, 8'd128, 8'd108, 8'd105, 8'd155, 8'd103, 8'd94, 8'd108, 8'd102, 8'd48, 8'd96, 8'd136, 8'd91, 8'd90, 8'd117, 8'd82, 8'd73, 8'd77, 8'd59, 8'd145, 8'd136, 8'd177, 8'd153, 8'd102, 8'd97, 8'd125, 8'd107, 8'd120, 8'd92, 8'd150, 8'd116, 8'd142, 8'd138, 8'd97, 8'd81, 8'd160, 8'd150, 8'd67, 8'd137, 8'd117, 8'd127, 8'd122, 8'd90, 8'd101, 8'd70, 8'd108, 8'd91, 8'd117, 8'd146, 8'd141, 8'd84, 8'd93, 8'd115, 8'd120, 8'd110, 8'd115, 8'd67, 8'd101, 8'd87, 8'd100, 8'd96, 8'd165, 8'd133, 8'd139, 8'd171, 8'd140, 8'd105, 8'd152, 8'd149, 8'd62, 8'd45, 8'd65, 8'd76, 8'd72, 8'd70, 8'd80, 8'd156, 8'd124, 8'd159, 8'd138, 8'd45, 8'd45, 8'd65, 8'd109, 8'd67, 8'd119, 8'd116, 8'd147, 8'd74, 8'd180, 8'd131, 8'd205, 8'd154, 8'd146, 8'd119, 8'd98, 8'd168, 8'd132, 8'd113, 8'd112, 8'd73, 8'd122, 8'd66, 8'd120, 8'd93, 8'd80, 8'd119, 8'd59, 8'd87, 8'd98, 8'd96, 8'd125, 8'd111, 8'd92, 8'd71, 8'd105, 8'd137, 8'd153, 8'd124, 8'd153, 8'd153, 8'd98, 8'd75, 8'd159, 8'd160, 8'd113, 8'd78, 8'd119, 8'd93, 8'd135, 8'd113, 8'd95, 8'd87, 8'd102, 8'd102, 8'd87, 8'd67, 8'd41, 8'd108, 8'd73, 8'd94, 8'd171, 8'd178, 8'd184, 8'd160, 8'd163, 8'd188, 8'd152, 8'd85, 8'd65, 8'd51, 8'd127, 8'd136, 8'd120, 8'd132, 8'd123, 8'd111, 8'd141, 8'd154, 8'd79, 8'd139, 8'd135, 8'd129, 8'd134, 8'd58, 8'd105, 8'd152, 8'd93, 8'd152, 8'd102, 8'd109, 8'd162, 8'd111, 8'd178, 8'd174, 8'd106, 8'd94, 8'd110, 8'd91, 8'd115, 8'd87, 8'd143, 8'd131, 8'd170, 8'd90, 8'd148, 8'd131, 8'd94, 8'd78, 8'd133, 8'd86, 8'd88, 8'd128, 8'd77, 8'd102, 8'd137, 8'd181, 8'd138, 8'd182, 8'd184, 8'd167, 8'd208, 8'd155, 8'd120, 8'd61, 8'd66, 8'd141, 8'd91, 8'd90, 8'd132, 8'd78, 8'd93, 8'd169, 8'd161, 8'd147, 8'd168, 8'd118, 8'd141, 8'd132, 8'd128, 8'd151, 8'd182, 8'd185, 8'd113, 8'd168, 8'd181, 8'd166, 8'd128, 8'd155, 8'd134, 8'd198, 8'd107, 8'd115, 8'd144, 8'd151, 8'd139, 8'd189, 8'd123, 8'd160, 8'd126, 8'd173, 8'd137, 8'd88, 8'd130, 8'd85, 8'd158, 8'd82, 8'd67, 8'd137, 8'd143, 8'd169, 8'd130, 8'd168, 8'd152, 8'd147, 8'd151, 8'd199, 8'd163, 8'd104, 8'd126, 8'd139, 8'd86, 8'd122, 8'd136, 8'd98, 8'd158, 8'd124, 8'd133, 8'd137, 8'd162, 8'd174, 8'd136, 8'd116, 8'd100, 8'd97, 8'd95, 8'd44, 8'd98, 8'd161, 8'd118, 8'd128, 8'd119, 8'd150, 8'd105, 8'd122, 8'd90, 8'd161, 8'd116, 8'd72, 8'd127, 8'd121, 8'd90, 8'd171, 8'd106, 8'd110, 8'd124, 8'd149, 8'd138, 8'd97, 8'd157, 8'd98, 8'd135, 8'd69, 8'd83, 8'd79, 8'd134, 8'd116, 8'd108, 8'd132, 8'd112, 8'd144, 8'd115, 8'd142, 8'd86, 8'd116, 8'd162, 8'd138, 8'd116, 8'd148, 8'd88, 8'd100, 8'd153, 8'd87, 8'd105, 8'd172, 8'd107, 8'd158, 8'd126, 8'd79, 8'd122, 8'd155, 8'd131, 8'd136, 8'd95, 8'd83, 8'd89, 8'd75, 8'd161, 8'd123, 8'd141, 8'd126, 8'd92, 8'd156, 8'd148, 8'd127, 8'd115, 8'd124, 8'd121, 8'd130, 8'd158, 8'd164, 8'd108, 8'd140, 8'd101, 8'd142, 8'd154, 8'd130, 8'd92, 8'd78, 8'd57, 8'd107, 8'd71, 8'd69, 8'd83, 8'd118, 8'd100, 8'd134, 8'd113, 8'd75, 8'd136, 8'd134, 8'd159, 8'd145, 8'd91, 8'd105, 8'd156, 8'd102, 8'd137, 8'd160, 8'd86, 8'd116, 8'd136, 8'd78, 8'd61, 8'd120, 8'd60, 8'd65, 8'd77, 8'd112, 8'd157, 8'd110, 8'd154, 8'd164, 8'd127, 8'd64, 8'd151, 8'd57, 8'd126, 8'd104, 8'd101, 8'd127, 8'd109, 8'd108, 8'd167, 8'd158, 8'd140, 8'd77, 8'd128, 8'd180, 8'd116, 8'd89, 8'd107, 8'd114, 8'd148, 8'd94, 8'd122, 8'd150, 8'd74, 8'd108, 8'd163, 8'd125, 8'd93, 8'd74, 8'd111, 8'd57, 8'd79, 8'd157, 8'd153, 8'd72, 8'd65, 8'd115, 8'd83, 8'd83, 8'd165, 8'd148, 8'd154, 8'd155, 8'd89, 8'd124, 8'd134, 8'd154, 8'd155, 8'd143, 8'd96, 8'd126, 8'd157, 8'd137, 8'd82, 8'd128, 8'd151, 8'd135, 8'd133, 8'd68, 8'd124, 8'd76, 8'd153, 8'd57, 8'd76, 8'd123, 8'd101, 8'd149, 8'd113, 8'd83, 8'd123, 8'd179, 8'd78, 8'd114, 8'd119, 8'd96, 8'd165, 8'd80, 8'd125, 8'd99, 8'd81, 8'd152, 8'd101, 8'd55, 8'd134, 8'd97, 8'd137, 8'd83, 8'd143, 8'd127, 8'd121, 8'd107, 8'd82, 8'd107, 8'd134, 8'd57, 8'd134, 8'd167, 8'd139, 8'd115, 8'd106, 8'd173, 8'd115, 8'd157, 8'd106, 8'd156, 8'd123, 8'd126, 8'd74, 8'd169, 8'd97, 8'd121, 8'd136, 8'd69, 8'd67, 8'd75, 8'd153, 8'd121, 8'd122, 8'd129, 8'd116, 8'd112, 8'd120, 8'd112, 8'd125, 8'd140, 8'd79, 8'd130, 8'd164, 8'd102, 8'd152, 8'd167, 8'd150, 8'd134, 8'd154, 8'd155, 8'd145, 8'd126, 8'd122, 8'd79, 8'd158, 8'd97, 8'd97, 8'd90, 8'd141, 8'd133, 8'd122, 8'd108, 8'd100, 8'd124, 8'd94, 8'd87, 8'd96, 8'd77, 8'd88, 8'd148, 8'd80, 8'd157, 8'd118, 8'd116, 8'd78, 8'd146, 8'd70, 8'd125, 8'd167, 8'd117, 8'd139, 8'd147, 8'd138, 8'd76, 8'd87, 8'd124, 8'd156, 8'd117, 8'd131, 8'd78, 8'd112, 8'd99, 8'd120, 8'd109, 8'd161, 8'd163, 8'd165, 8'd153, 8'd75, 8'd101, 8'd100, 8'd142})
) cell_0_10 (
    .clk(clk),
    .input_index(index_0_9_10),
    .input_value(value_0_9_10),
    .input_result(result_0_9_10),
    .input_enable(enable_0_9_10),
    .output_index(index_0_10_11),
    .output_value(value_0_10_11),
    .output_result(result_0_10_11),
    .output_enable(enable_0_10_11)
);

wire [10-1:0] index_0_11_12;
wire [`DATA_WIDTH-1:0] value_0_11_12;
wire [`DATA_WIDTH*4:0] result_0_11_12;
wire enable_0_11_12;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd89, 8'd122, 8'd71, 8'd78, 8'd148, 8'd162, 8'd155, 8'd127, 8'd155, 8'd116, 8'd196, 8'd158, 8'd139, 8'd201, 8'd191, 8'd129, 8'd106, 8'd131, 8'd106, 8'd132, 8'd86, 8'd131, 8'd157, 8'd124, 8'd118, 8'd167, 8'd76, 8'd120, 8'd124, 8'd140, 8'd143, 8'd157, 8'd152, 8'd188, 8'd189, 8'd137, 8'd209, 8'd158, 8'd193, 8'd175, 8'd142, 8'd229, 8'd154, 8'd201, 8'd191, 8'd196, 8'd200, 8'd205, 8'd148, 8'd141, 8'd108, 8'd91, 8'd168, 8'd166, 8'd158, 8'd158, 8'd138, 8'd161, 8'd143, 8'd95, 8'd136, 8'd174, 8'd186, 8'd123, 8'd128, 8'd200, 8'd228, 8'd181, 8'd168, 8'd176, 8'd209, 8'd206, 8'd221, 8'd227, 8'd161, 8'd167, 8'd138, 8'd134, 8'd103, 8'd138, 8'd94, 8'd158, 8'd148, 8'd158, 8'd105, 8'd102, 8'd124, 8'd70, 8'd98, 8'd122, 8'd184, 8'd199, 8'd154, 8'd176, 8'd106, 8'd187, 8'd150, 8'd166, 8'd177, 8'd188, 8'd126, 8'd134, 8'd120, 8'd177, 8'd111, 8'd161, 8'd164, 8'd141, 8'd124, 8'd119, 8'd157, 8'd104, 8'd77, 8'd94, 8'd120, 8'd111, 8'd79, 8'd140, 8'd162, 8'd89, 8'd179, 8'd162, 8'd106, 8'd192, 8'd177, 8'd161, 8'd166, 8'd143, 8'd99, 8'd79, 8'd137, 8'd82, 8'd80, 8'd98, 8'd111, 8'd126, 8'd70, 8'd71, 8'd139, 8'd109, 8'd67, 8'd81, 8'd143, 8'd118, 8'd82, 8'd150, 8'd158, 8'd139, 8'd108, 8'd126, 8'd114, 8'd113, 8'd137, 8'd89, 8'd140, 8'd119, 8'd84, 8'd152, 8'd118, 8'd135, 8'd140, 8'd102, 8'd92, 8'd85, 8'd89, 8'd145, 8'd95, 8'd85, 8'd90, 8'd136, 8'd77, 8'd149, 8'd117, 8'd105, 8'd153, 8'd120, 8'd91, 8'd87, 8'd131, 8'd76, 8'd89, 8'd93, 8'd60, 8'd50, 8'd75, 8'd94, 8'd67, 8'd70, 8'd148, 8'd148, 8'd149, 8'd92, 8'd96, 8'd99, 8'd75, 8'd99, 8'd171, 8'd94, 8'd138, 8'd120, 8'd157, 8'd128, 8'd67, 8'd64, 8'd92, 8'd135, 8'd100, 8'd127, 8'd123, 8'd102, 8'd98, 8'd55, 8'd101, 8'd110, 8'd103, 8'd116, 8'd150, 8'd162, 8'd146, 8'd141, 8'd140, 8'd159, 8'd99, 8'd110, 8'd127, 8'd97, 8'd79, 8'd150, 8'd74, 8'd124, 8'd93, 8'd117, 8'd128, 8'd147, 8'd149, 8'd136, 8'd137, 8'd99, 8'd82, 8'd43, 8'd87, 8'd106, 8'd63, 8'd84, 8'd70, 8'd126, 8'd163, 8'd74, 8'd160, 8'd174, 8'd101, 8'd132, 8'd134, 8'd69, 8'd115, 8'd92, 8'd67, 8'd146, 8'd136, 8'd113, 8'd142, 8'd73, 8'd156, 8'd115, 8'd159, 8'd117, 8'd151, 8'd63, 8'd60, 8'd36, 8'd98, 8'd148, 8'd148, 8'd152, 8'd66, 8'd140, 8'd126, 8'd100, 8'd172, 8'd99, 8'd128, 8'd89, 8'd57, 8'd62, 8'd64, 8'd80, 8'd103, 8'd128, 8'd106, 8'd136, 8'd173, 8'd176, 8'd183, 8'd150, 8'd157, 8'd86, 8'd104, 8'd70, 8'd43, 8'd127, 8'd114, 8'd116, 8'd143, 8'd121, 8'd115, 8'd169, 8'd158, 8'd117, 8'd74, 8'd42, 8'd37, 8'd118, 8'd130, 8'd114, 8'd112, 8'd149, 8'd147, 8'd140, 8'd122, 8'd194, 8'd183, 8'd121, 8'd196, 8'd111, 8'd88, 8'd89, 8'd88, 8'd125, 8'd71, 8'd88, 8'd96, 8'd89, 8'd103, 8'd124, 8'd154, 8'd138, 8'd126, 8'd97, 8'd113, 8'd118, 8'd109, 8'd101, 8'd104, 8'd133, 8'd126, 8'd168, 8'd109, 8'd198, 8'd119, 8'd205, 8'd153, 8'd123, 8'd104, 8'd105, 8'd90, 8'd66, 8'd38, 8'd80, 8'd95, 8'd118, 8'd141, 8'd107, 8'd96, 8'd97, 8'd144, 8'd126, 8'd65, 8'd71, 8'd77, 8'd58, 8'd148, 8'd98, 8'd145, 8'd183, 8'd114, 8'd167, 8'd194, 8'd163, 8'd128, 8'd151, 8'd75, 8'd28, 8'd120, 8'd58, 8'd67, 8'd71, 8'd135, 8'd179, 8'd158, 8'd175, 8'd159, 8'd110, 8'd79, 8'd95, 8'd109, 8'd29, 8'd108, 8'd110, 8'd72, 8'd106, 8'd118, 8'd166, 8'd133, 8'd213, 8'd153, 8'd142, 8'd176, 8'd150, 8'd127, 8'd86, 8'd109, 8'd92, 8'd166, 8'd133, 8'd185, 8'd201, 8'd129, 8'd94, 8'd96, 8'd149, 8'd104, 8'd181, 8'd164, 8'd114, 8'd74, 8'd97, 8'd106, 8'd90, 8'd116, 8'd158, 8'd165, 8'd168, 8'd222, 8'd217, 8'd115, 8'd130, 8'd141, 8'd142, 8'd153, 8'd123, 8'd162, 8'd176, 8'd117, 8'd122, 8'd121, 8'd172, 8'd160, 8'd152, 8'd107, 8'd198, 8'd132, 8'd147, 8'd73, 8'd113, 8'd129, 8'd76, 8'd131, 8'd194, 8'd172, 8'd154, 8'd173, 8'd191, 8'd108, 8'd139, 8'd166, 8'd154, 8'd137, 8'd164, 8'd165, 8'd144, 8'd200, 8'd201, 8'd135, 8'd165, 8'd113, 8'd142, 8'd125, 8'd163, 8'd181, 8'd77, 8'd137, 8'd149, 8'd102, 8'd160, 8'd105, 8'd146, 8'd130, 8'd117, 8'd177, 8'd170, 8'd83, 8'd114, 8'd126, 8'd107, 8'd194, 8'd110, 8'd137, 8'd173, 8'd159, 8'd194, 8'd86, 8'd160, 8'd169, 8'd79, 8'd153, 8'd184, 8'd210, 8'd156, 8'd103, 8'd103, 8'd182, 8'd130, 8'd132, 8'd158, 8'd121, 8'd97, 8'd131, 8'd94, 8'd144, 8'd131, 8'd147, 8'd121, 8'd195, 8'd110, 8'd110, 8'd187, 8'd127, 8'd132, 8'd96, 8'd85, 8'd155, 8'd159, 8'd123, 8'd163, 8'd223, 8'd177, 8'd98, 8'd113, 8'd122, 8'd137, 8'd154, 8'd184, 8'd115, 8'd118, 8'd141, 8'd114, 8'd126, 8'd149, 8'd108, 8'd144, 8'd170, 8'd183, 8'd115, 8'd183, 8'd181, 8'd129, 8'd165, 8'd79, 8'd78, 8'd148, 8'd163, 8'd103, 8'd168, 8'd100, 8'd107, 8'd159, 8'd165, 8'd96, 8'd146, 8'd137, 8'd120, 8'd113, 8'd146, 8'd102, 8'd148, 8'd147, 8'd189, 8'd151, 8'd152, 8'd114, 8'd102, 8'd157, 8'd74, 8'd76, 8'd107, 8'd112, 8'd92, 8'd80, 8'd100, 8'd176, 8'd202, 8'd154, 8'd140, 8'd114, 8'd106, 8'd161, 8'd102, 8'd82, 8'd146, 8'd113, 8'd143, 8'd123, 8'd80, 8'd88, 8'd148, 8'd162, 8'd86, 8'd141, 8'd85, 8'd114, 8'd120, 8'd122, 8'd90, 8'd174, 8'd150, 8'd79, 8'd112, 8'd167, 8'd119, 8'd174, 8'd150, 8'd99, 8'd91, 8'd113, 8'd61, 8'd56, 8'd52, 8'd114, 8'd98, 8'd142, 8'd68, 8'd110, 8'd103, 8'd164, 8'd146, 8'd143, 8'd134, 8'd133, 8'd117, 8'd74, 8'd120, 8'd123, 8'd109, 8'd156, 8'd119, 8'd165, 8'd150, 8'd78, 8'd147, 8'd97, 8'd128, 8'd75, 8'd86, 8'd106, 8'd72, 8'd128, 8'd86, 8'd144, 8'd84, 8'd84, 8'd127, 8'd136, 8'd91, 8'd61, 8'd117, 8'd151, 8'd87, 8'd118, 8'd163, 8'd138, 8'd89, 8'd123, 8'd163, 8'd118, 8'd74, 8'd71, 8'd101, 8'd151, 8'd79, 8'd74, 8'd147, 8'd154, 8'd73, 8'd94, 8'd100, 8'd97, 8'd60, 8'd106, 8'd77, 8'd50, 8'd55, 8'd79, 8'd102, 8'd125, 8'd93, 8'd76, 8'd144, 8'd101, 8'd115, 8'd75, 8'd82, 8'd164, 8'd96, 8'd83, 8'd133, 8'd109, 8'd130, 8'd87, 8'd104, 8'd74, 8'd84, 8'd118, 8'd79, 8'd112, 8'd99, 8'd91, 8'd46, 8'd67, 8'd79, 8'd53, 8'd139, 8'd97, 8'd74, 8'd87, 8'd160, 8'd156, 8'd137, 8'd148, 8'd112, 8'd76, 8'd94, 8'd154, 8'd106, 8'd93, 8'd119, 8'd101, 8'd141, 8'd108, 8'd92, 8'd112, 8'd108, 8'd73, 8'd133, 8'd50, 8'd51, 8'd126, 8'd97, 8'd150, 8'd145, 8'd70, 8'd116, 8'd76, 8'd167, 8'd168, 8'd84, 8'd70, 8'd167, 8'd117, 8'd80, 8'd98, 8'd110, 8'd94, 8'd167, 8'd166, 8'd104, 8'd75, 8'd72, 8'd137, 8'd94, 8'd128, 8'd111, 8'd119, 8'd78, 8'd130, 8'd139, 8'd126, 8'd158, 8'd115, 8'd117, 8'd88, 8'd74, 8'd161, 8'd153, 8'd91})
) cell_0_11 (
    .clk(clk),
    .input_index(index_0_10_11),
    .input_value(value_0_10_11),
    .input_result(result_0_10_11),
    .input_enable(enable_0_10_11),
    .output_index(index_0_11_12),
    .output_value(value_0_11_12),
    .output_result(result_0_11_12),
    .output_enable(enable_0_11_12)
);

wire [10-1:0] index_0_12_13;
wire [`DATA_WIDTH-1:0] value_0_12_13;
wire [`DATA_WIDTH*4:0] result_0_12_13;
wire enable_0_12_13;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd108, 8'd105, 8'd145, 8'd100, 8'd83, 8'd113, 8'd88, 8'd77, 8'd78, 8'd97, 8'd67, 8'd101, 8'd146, 8'd139, 8'd127, 8'd60, 8'd140, 8'd94, 8'd130, 8'd67, 8'd160, 8'd78, 8'd144, 8'd83, 8'd135, 8'd100, 8'd102, 8'd94, 8'd119, 8'd98, 8'd97, 8'd145, 8'd140, 8'd70, 8'd100, 8'd117, 8'd132, 8'd102, 8'd113, 8'd139, 8'd58, 8'd145, 8'd104, 8'd73, 8'd62, 8'd123, 8'd101, 8'd122, 8'd135, 8'd79, 8'd112, 8'd107, 8'd150, 8'd169, 8'd157, 8'd92, 8'd93, 8'd130, 8'd171, 8'd130, 8'd158, 8'd148, 8'd162, 8'd102, 8'd78, 8'd118, 8'd70, 8'd86, 8'd113, 8'd85, 8'd87, 8'd81, 8'd80, 8'd62, 8'd51, 8'd106, 8'd93, 8'd126, 8'd128, 8'd115, 8'd64, 8'd122, 8'd136, 8'd148, 8'd130, 8'd150, 8'd118, 8'd85, 8'd107, 8'd144, 8'd112, 8'd147, 8'd102, 8'd163, 8'd88, 8'd95, 8'd112, 8'd75, 8'd91, 8'd66, 8'd132, 8'd116, 8'd110, 8'd61, 8'd115, 8'd49, 8'd51, 8'd86, 8'd103, 8'd122, 8'd155, 8'd122, 8'd110, 8'd113, 8'd131, 8'd145, 8'd121, 8'd179, 8'd161, 8'd135, 8'd146, 8'd102, 8'd141, 8'd146, 8'd120, 8'd132, 8'd98, 8'd81, 8'd75, 8'd90, 8'd98, 8'd117, 8'd96, 8'd84, 8'd143, 8'd87, 8'd119, 8'd102, 8'd116, 8'd142, 8'd166, 8'd72, 8'd98, 8'd151, 8'd116, 8'd121, 8'd129, 8'd151, 8'd127, 8'd152, 8'd97, 8'd148, 8'd104, 8'd78, 8'd106, 8'd129, 8'd112, 8'd105, 8'd139, 8'd90, 8'd131, 8'd137, 8'd101, 8'd85, 8'd167, 8'd140, 8'd77, 8'd111, 8'd128, 8'd143, 8'd103, 8'd95, 8'd117, 8'd102, 8'd115, 8'd175, 8'd107, 8'd96, 8'd140, 8'd127, 8'd90, 8'd162, 8'd155, 8'd97, 8'd95, 8'd144, 8'd95, 8'd151, 8'd168, 8'd125, 8'd144, 8'd156, 8'd147, 8'd88, 8'd76, 8'd110, 8'd158, 8'd167, 8'd164, 8'd158, 8'd159, 8'd141, 8'd104, 8'd136, 8'd152, 8'd136, 8'd83, 8'd113, 8'd143, 8'd96, 8'd158, 8'd127, 8'd138, 8'd108, 8'd130, 8'd168, 8'd138, 8'd164, 8'd84, 8'd104, 8'd120, 8'd104, 8'd147, 8'd160, 8'd153, 8'd100, 8'd184, 8'd93, 8'd101, 8'd95, 8'd125, 8'd116, 8'd153, 8'd93, 8'd178, 8'd108, 8'd112, 8'd95, 8'd135, 8'd127, 8'd107, 8'd132, 8'd118, 8'd178, 8'd100, 8'd123, 8'd144, 8'd142, 8'd130, 8'd148, 8'd85, 8'd126, 8'd131, 8'd151, 8'd183, 8'd197, 8'd94, 8'd135, 8'd104, 8'd101, 8'd108, 8'd173, 8'd136, 8'd93, 8'd102, 8'd156, 8'd149, 8'd160, 8'd116, 8'd109, 8'd165, 8'd118, 8'd172, 8'd94, 8'd108, 8'd128, 8'd132, 8'd97, 8'd151, 8'd108, 8'd188, 8'd171, 8'd214, 8'd107, 8'd102, 8'd87, 8'd100, 8'd122, 8'd152, 8'd77, 8'd73, 8'd84, 8'd101, 8'd106, 8'd130, 8'd172, 8'd107, 8'd158, 8'd128, 8'd135, 8'd167, 8'd116, 8'd91, 8'd140, 8'd166, 8'd129, 8'd107, 8'd146, 8'd155, 8'd120, 8'd147, 8'd145, 8'd148, 8'd105, 8'd117, 8'd157, 8'd98, 8'd101, 8'd160, 8'd177, 8'd158, 8'd182, 8'd145, 8'd149, 8'd176, 8'd187, 8'd94, 8'd118, 8'd129, 8'd163, 8'd86, 8'd139, 8'd134, 8'd81, 8'd129, 8'd140, 8'd180, 8'd166, 8'd171, 8'd104, 8'd155, 8'd57, 8'd73, 8'd114, 8'd63, 8'd58, 8'd161, 8'd112, 8'd124, 8'd164, 8'd152, 8'd117, 8'd126, 8'd154, 8'd95, 8'd124, 8'd109, 8'd93, 8'd88, 8'd81, 8'd159, 8'd151, 8'd95, 8'd67, 8'd145, 8'd137, 8'd148, 8'd102, 8'd148, 8'd103, 8'd87, 8'd142, 8'd111, 8'd86, 8'd81, 8'd172, 8'd87, 8'd176, 8'd132, 8'd157, 8'd166, 8'd88, 8'd97, 8'd132, 8'd135, 8'd100, 8'd132, 8'd90, 8'd127, 8'd85, 8'd111, 8'd99, 8'd107, 8'd143, 8'd128, 8'd124, 8'd202, 8'd120, 8'd129, 8'd113, 8'd132, 8'd169, 8'd78, 8'd83, 8'd128, 8'd164, 8'd137, 8'd80, 8'd85, 8'd149, 8'd60, 8'd100, 8'd123, 8'd128, 8'd120, 8'd120, 8'd76, 8'd119, 8'd81, 8'd121, 8'd174, 8'd89, 8'd87, 8'd226, 8'd146, 8'd148, 8'd153, 8'd109, 8'd173, 8'd125, 8'd132, 8'd83, 8'd150, 8'd117, 8'd90, 8'd98, 8'd141, 8'd79, 8'd71, 8'd81, 8'd75, 8'd99, 8'd120, 8'd139, 8'd102, 8'd48, 8'd77, 8'd145, 8'd68, 8'd71, 8'd119, 8'd72, 8'd113, 8'd125, 8'd108, 8'd109, 8'd136, 8'd149, 8'd88, 8'd96, 8'd102, 8'd135, 8'd97, 8'd135, 8'd57, 8'd64, 8'd91, 8'd135, 8'd93, 8'd95, 8'd162, 8'd76, 8'd71, 8'd48, 8'd53, 8'd118, 8'd125, 8'd129, 8'd93, 8'd102, 8'd148, 8'd100, 8'd99, 8'd99, 8'd155, 8'd85, 8'd80, 8'd69, 8'd145, 8'd74, 8'd116, 8'd78, 8'd121, 8'd116, 8'd108, 8'd108, 8'd96, 8'd137, 8'd123, 8'd153, 8'd150, 8'd134, 8'd151, 8'd103, 8'd96, 8'd100, 8'd120, 8'd52, 8'd96, 8'd109, 8'd156, 8'd107, 8'd105, 8'd98, 8'd135, 8'd126, 8'd120, 8'd115, 8'd113, 8'd80, 8'd109, 8'd110, 8'd124, 8'd111, 8'd117, 8'd119, 8'd154, 8'd159, 8'd87, 8'd85, 8'd145, 8'd131, 8'd90, 8'd139, 8'd59, 8'd89, 8'd60, 8'd110, 8'd137, 8'd146, 8'd98, 8'd128, 8'd147, 8'd108, 8'd103, 8'd83, 8'd125, 8'd87, 8'd152, 8'd76, 8'd76, 8'd139, 8'd81, 8'd171, 8'd128, 8'd90, 8'd153, 8'd141, 8'd150, 8'd106, 8'd80, 8'd131, 8'd113, 8'd91, 8'd116, 8'd135, 8'd144, 8'd102, 8'd116, 8'd157, 8'd107, 8'd130, 8'd172, 8'd181, 8'd120, 8'd151, 8'd122, 8'd161, 8'd89, 8'd137, 8'd122, 8'd89, 8'd94, 8'd172, 8'd105, 8'd137, 8'd75, 8'd157, 8'd114, 8'd111, 8'd128, 8'd64, 8'd115, 8'd67, 8'd77, 8'd139, 8'd157, 8'd120, 8'd155, 8'd163, 8'd129, 8'd175, 8'd151, 8'd78, 8'd169, 8'd116, 8'd91, 8'd93, 8'd151, 8'd140, 8'd92, 8'd109, 8'd136, 8'd145, 8'd161, 8'd83, 8'd90, 8'd86, 8'd92, 8'd88, 8'd118, 8'd122, 8'd151, 8'd79, 8'd134, 8'd107, 8'd140, 8'd117, 8'd143, 8'd96, 8'd147, 8'd132, 8'd113, 8'd184, 8'd157, 8'd126, 8'd136, 8'd133, 8'd163, 8'd129, 8'd144, 8'd132, 8'd129, 8'd141, 8'd130, 8'd91, 8'd128, 8'd88, 8'd100, 8'd53, 8'd79, 8'd69, 8'd144, 8'd94, 8'd89, 8'd143, 8'd96, 8'd161, 8'd182, 8'd125, 8'd156, 8'd174, 8'd149, 8'd158, 8'd132, 8'd99, 8'd149, 8'd123, 8'd68, 8'd123, 8'd101, 8'd72, 8'd157, 8'd163, 8'd101, 8'd137, 8'd161, 8'd79, 8'd142, 8'd108, 8'd123, 8'd106, 8'd115, 8'd152, 8'd156, 8'd103, 8'd124, 8'd138, 8'd145, 8'd166, 8'd161, 8'd180, 8'd145, 8'd165, 8'd156, 8'd76, 8'd110, 8'd136, 8'd79, 8'd110, 8'd156, 8'd83, 8'd164, 8'd111, 8'd119, 8'd137, 8'd146, 8'd128, 8'd90, 8'd178, 8'd169, 8'd128, 8'd132, 8'd182, 8'd192, 8'd148, 8'd201, 8'd147, 8'd116, 8'd192, 8'd144, 8'd105, 8'd126, 8'd150, 8'd176, 8'd153, 8'd76, 8'd134, 8'd78, 8'd166, 8'd83, 8'd126, 8'd87, 8'd101, 8'd169, 8'd142, 8'd177, 8'd157, 8'd101, 8'd140, 8'd126, 8'd138, 8'd155, 8'd130, 8'd166, 8'd121, 8'd85, 8'd99, 8'd143, 8'd154, 8'd159, 8'd107, 8'd154, 8'd86, 8'd136, 8'd95, 8'd116, 8'd127, 8'd121, 8'd120, 8'd87, 8'd101, 8'd145, 8'd72, 8'd84, 8'd72, 8'd164, 8'd160, 8'd159, 8'd155, 8'd92, 8'd149, 8'd86, 8'd103, 8'd155, 8'd77, 8'd153, 8'd155, 8'd75, 8'd161, 8'd92, 8'd155, 8'd118, 8'd87})
) cell_0_12 (
    .clk(clk),
    .input_index(index_0_11_12),
    .input_value(value_0_11_12),
    .input_result(result_0_11_12),
    .input_enable(enable_0_11_12),
    .output_index(index_0_12_13),
    .output_value(value_0_12_13),
    .output_result(result_0_12_13),
    .output_enable(enable_0_12_13)
);

wire [10-1:0] index_0_13_14;
wire [`DATA_WIDTH-1:0] value_0_13_14;
wire [`DATA_WIDTH*4:0] result_0_13_14;
wire enable_0_13_14;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd82, 8'd147, 8'd136, 8'd95, 8'd162, 8'd104, 8'd150, 8'd129, 8'd183, 8'd103, 8'd154, 8'd173, 8'd141, 8'd102, 8'd175, 8'd176, 8'd146, 8'd106, 8'd130, 8'd89, 8'd131, 8'd165, 8'd146, 8'd157, 8'd123, 8'd130, 8'd157, 8'd106, 8'd101, 8'd161, 8'd126, 8'd82, 8'd116, 8'd132, 8'd84, 8'd174, 8'd163, 8'd142, 8'd167, 8'd166, 8'd117, 8'd121, 8'd188, 8'd179, 8'd165, 8'd90, 8'd149, 8'd169, 8'd106, 8'd112, 8'd118, 8'd120, 8'd94, 8'd143, 8'd169, 8'd137, 8'd111, 8'd92, 8'd61, 8'd109, 8'd171, 8'd116, 8'd100, 8'd137, 8'd131, 8'd190, 8'd126, 8'd124, 8'd123, 8'd132, 8'd126, 8'd206, 8'd190, 8'd126, 8'd122, 8'd187, 8'd160, 8'd182, 8'd119, 8'd138, 8'd121, 8'd119, 8'd71, 8'd142, 8'd148, 8'd107, 8'd112, 8'd97, 8'd53, 8'd97, 8'd76, 8'd168, 8'd166, 8'd116, 8'd113, 8'd153, 8'd193, 8'd194, 8'd141, 8'd122, 8'd134, 8'd192, 8'd115, 8'd136, 8'd136, 8'd120, 8'd127, 8'd178, 8'd130, 8'd147, 8'd116, 8'd119, 8'd130, 8'd113, 8'd63, 8'd110, 8'd49, 8'd93, 8'd102, 8'd92, 8'd106, 8'd171, 8'd185, 8'd130, 8'd90, 8'd148, 8'd162, 8'd133, 8'd150, 8'd86, 8'd77, 8'd75, 8'd169, 8'd162, 8'd133, 8'd156, 8'd119, 8'd82, 8'd126, 8'd78, 8'd163, 8'd130, 8'd105, 8'd59, 8'd54, 8'd45, 8'd154, 8'd115, 8'd137, 8'd148, 8'd79, 8'd149, 8'd168, 8'd140, 8'd118, 8'd79, 8'd103, 8'd150, 8'd96, 8'd148, 8'd81, 8'd115, 8'd94, 8'd101, 8'd110, 8'd130, 8'd119, 8'd125, 8'd114, 8'd77, 8'd139, 8'd130, 8'd107, 8'd84, 8'd129, 8'd124, 8'd145, 8'd160, 8'd136, 8'd102, 8'd103, 8'd101, 8'd153, 8'd88, 8'd94, 8'd149, 8'd85, 8'd157, 8'd85, 8'd74, 8'd74, 8'd63, 8'd101, 8'd121, 8'd121, 8'd164, 8'd133, 8'd102, 8'd116, 8'd145, 8'd109, 8'd149, 8'd135, 8'd95, 8'd159, 8'd90, 8'd137, 8'd108, 8'd96, 8'd139, 8'd154, 8'd136, 8'd69, 8'd147, 8'd61, 8'd100, 8'd114, 8'd103, 8'd104, 8'd62, 8'd99, 8'd119, 8'd125, 8'd103, 8'd174, 8'd65, 8'd139, 8'd135, 8'd61, 8'd107, 8'd99, 8'd144, 8'd137, 8'd138, 8'd97, 8'd108, 8'd82, 8'd133, 8'd88, 8'd158, 8'd126, 8'd53, 8'd123, 8'd92, 8'd111, 8'd79, 8'd66, 8'd125, 8'd170, 8'd106, 8'd103, 8'd122, 8'd152, 8'd108, 8'd51, 8'd89, 8'd119, 8'd65, 8'd84, 8'd133, 8'd131, 8'd91, 8'd75, 8'd153, 8'd97, 8'd116, 8'd102, 8'd135, 8'd77, 8'd108, 8'd69, 8'd87, 8'd79, 8'd118, 8'd67, 8'd148, 8'd101, 8'd163, 8'd97, 8'd114, 8'd146, 8'd65, 8'd38, 8'd71, 8'd105, 8'd95, 8'd131, 8'd138, 8'd125, 8'd86, 8'd123, 8'd90, 8'd141, 8'd102, 8'd138, 8'd144, 8'd55, 8'd124, 8'd126, 8'd116, 8'd50, 8'd101, 8'd71, 8'd89, 8'd172, 8'd157, 8'd176, 8'd168, 8'd124, 8'd97, 8'd74, 8'd94, 8'd75, 8'd103, 8'd155, 8'd149, 8'd139, 8'd99, 8'd151, 8'd185, 8'd110, 8'd132, 8'd114, 8'd149, 8'd66, 8'd26, 8'd121, 8'd104, 8'd74, 8'd136, 8'd117, 8'd84, 8'd172, 8'd128, 8'd157, 8'd142, 8'd126, 8'd121, 8'd125, 8'd67, 8'd87, 8'd117, 8'd77, 8'd140, 8'd126, 8'd117, 8'd138, 8'd141, 8'd124, 8'd159, 8'd168, 8'd74, 8'd104, 8'd122, 8'd60, 8'd77, 8'd99, 8'd83, 8'd130, 8'd169, 8'd160, 8'd93, 8'd89, 8'd147, 8'd147, 8'd49, 8'd145, 8'd81, 8'd109, 8'd89, 8'd122, 8'd159, 8'd103, 8'd120, 8'd166, 8'd159, 8'd163, 8'd111, 8'd138, 8'd47, 8'd62, 8'd63, 8'd94, 8'd113, 8'd145, 8'd71, 8'd162, 8'd95, 8'd156, 8'd154, 8'd121, 8'd126, 8'd82, 8'd82, 8'd70, 8'd141, 8'd93, 8'd72, 8'd120, 8'd137, 8'd111, 8'd172, 8'd195, 8'd116, 8'd117, 8'd107, 8'd108, 8'd129, 8'd100, 8'd133, 8'd80, 8'd113, 8'd92, 8'd86, 8'd131, 8'd174, 8'd146, 8'd178, 8'd127, 8'd101, 8'd141, 8'd124, 8'd101, 8'd51, 8'd103, 8'd79, 8'd93, 8'd97, 8'd95, 8'd184, 8'd172, 8'd176, 8'd127, 8'd154, 8'd92, 8'd115, 8'd154, 8'd78, 8'd153, 8'd98, 8'd122, 8'd92, 8'd89, 8'd125, 8'd159, 8'd195, 8'd175, 8'd148, 8'd168, 8'd122, 8'd155, 8'd64, 8'd116, 8'd142, 8'd151, 8'd155, 8'd144, 8'd150, 8'd164, 8'd115, 8'd186, 8'd194, 8'd149, 8'd93, 8'd103, 8'd109, 8'd144, 8'd174, 8'd184, 8'd88, 8'd173, 8'd141, 8'd180, 8'd108, 8'd163, 8'd103, 8'd160, 8'd155, 8'd171, 8'd85, 8'd114, 8'd150, 8'd106, 8'd170, 8'd141, 8'd171, 8'd126, 8'd187, 8'd109, 8'd115, 8'd176, 8'd114, 8'd177, 8'd185, 8'd120, 8'd155, 8'd138, 8'd138, 8'd126, 8'd111, 8'd164, 8'd142, 8'd121, 8'd100, 8'd174, 8'd185, 8'd228, 8'd101, 8'd137, 8'd122, 8'd114, 8'd149, 8'd117, 8'd111, 8'd89, 8'd163, 8'd156, 8'd115, 8'd165, 8'd91, 8'd123, 8'd159, 8'd149, 8'd120, 8'd130, 8'd125, 8'd163, 8'd188, 8'd142, 8'd146, 8'd168, 8'd139, 8'd96, 8'd171, 8'd221, 8'd154, 8'd171, 8'd121, 8'd147, 8'd91, 8'd159, 8'd89, 8'd107, 8'd126, 8'd154, 8'd81, 8'd137, 8'd156, 8'd134, 8'd144, 8'd195, 8'd117, 8'd148, 8'd124, 8'd95, 8'd95, 8'd134, 8'd134, 8'd155, 8'd119, 8'd162, 8'd127, 8'd130, 8'd162, 8'd131, 8'd146, 8'd140, 8'd135, 8'd75, 8'd132, 8'd82, 8'd84, 8'd113, 8'd145, 8'd96, 8'd182, 8'd143, 8'd153, 8'd110, 8'd186, 8'd201, 8'd193, 8'd158, 8'd137, 8'd195, 8'd162, 8'd157, 8'd143, 8'd160, 8'd161, 8'd119, 8'd152, 8'd163, 8'd141, 8'd93, 8'd114, 8'd90, 8'd95, 8'd86, 8'd85, 8'd70, 8'd159, 8'd156, 8'd99, 8'd103, 8'd141, 8'd119, 8'd202, 8'd155, 8'd176, 8'd182, 8'd98, 8'd177, 8'd129, 8'd94, 8'd102, 8'd150, 8'd106, 8'd191, 8'd192, 8'd86, 8'd120, 8'd108, 8'd112, 8'd117, 8'd115, 8'd61, 8'd63, 8'd79, 8'd114, 8'd100, 8'd132, 8'd163, 8'd135, 8'd128, 8'd115, 8'd172, 8'd151, 8'd128, 8'd117, 8'd143, 8'd126, 8'd157, 8'd76, 8'd118, 8'd155, 8'd161, 8'd178, 8'd129, 8'd104, 8'd123, 8'd88, 8'd79, 8'd133, 8'd131, 8'd134, 8'd155, 8'd96, 8'd82, 8'd122, 8'd134, 8'd92, 8'd67, 8'd145, 8'd120, 8'd97, 8'd172, 8'd117, 8'd111, 8'd146, 8'd170, 8'd159, 8'd105, 8'd107, 8'd170, 8'd88, 8'd140, 8'd168, 8'd136, 8'd101, 8'd139, 8'd172, 8'd163, 8'd90, 8'd83, 8'd85, 8'd86, 8'd80, 8'd131, 8'd95, 8'd111, 8'd153, 8'd129, 8'd121, 8'd99, 8'd104, 8'd120, 8'd112, 8'd128, 8'd141, 8'd70, 8'd123, 8'd138, 8'd146, 8'd141, 8'd162, 8'd87, 8'd165, 8'd158, 8'd163, 8'd143, 8'd133, 8'd174, 8'd88, 8'd85, 8'd93, 8'd138, 8'd79, 8'd154, 8'd74, 8'd78, 8'd80, 8'd108, 8'd80, 8'd147, 8'd160, 8'd146, 8'd129, 8'd75, 8'd131, 8'd72, 8'd158, 8'd68, 8'd134, 8'd153, 8'd105, 8'd85, 8'd139, 8'd94, 8'd83, 8'd156, 8'd92, 8'd74, 8'd71, 8'd121, 8'd91, 8'd138, 8'd102, 8'd105, 8'd74, 8'd112, 8'd167, 8'd102, 8'd105, 8'd164, 8'd161, 8'd97, 8'd114, 8'd89, 8'd133, 8'd119, 8'd107, 8'd151, 8'd115, 8'd167, 8'd114, 8'd134, 8'd164, 8'd78, 8'd86, 8'd144, 8'd95, 8'd160, 8'd82, 8'd75, 8'd137, 8'd144, 8'd87, 8'd118, 8'd124, 8'd139, 8'd156, 8'd73, 8'd118})
) cell_0_13 (
    .clk(clk),
    .input_index(index_0_12_13),
    .input_value(value_0_12_13),
    .input_result(result_0_12_13),
    .input_enable(enable_0_12_13),
    .output_index(index_0_13_14),
    .output_value(value_0_13_14),
    .output_result(result_0_13_14),
    .output_enable(enable_0_13_14)
);

wire [10-1:0] index_0_14_15;
wire [`DATA_WIDTH-1:0] value_0_14_15;
wire [`DATA_WIDTH*4:0] result_0_14_15;
wire enable_0_14_15;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd141, 8'd90, 8'd98, 8'd118, 8'd142, 8'd169, 8'd127, 8'd117, 8'd130, 8'd137, 8'd164, 8'd164, 8'd137, 8'd179, 8'd119, 8'd120, 8'd131, 8'd147, 8'd109, 8'd169, 8'd92, 8'd128, 8'd75, 8'd109, 8'd113, 8'd158, 8'd70, 8'd111, 8'd135, 8'd83, 8'd146, 8'd82, 8'd162, 8'd155, 8'd107, 8'd131, 8'd143, 8'd111, 8'd161, 8'd168, 8'd212, 8'd183, 8'd164, 8'd174, 8'd213, 8'd145, 8'd145, 8'd159, 8'd165, 8'd149, 8'd182, 8'd99, 8'd88, 8'd160, 8'd91, 8'd153, 8'd74, 8'd119, 8'd113, 8'd154, 8'd88, 8'd160, 8'd103, 8'd121, 8'd119, 8'd189, 8'd159, 8'd162, 8'd126, 8'd168, 8'd177, 8'd132, 8'd130, 8'd143, 8'd168, 8'd187, 8'd130, 8'd185, 8'd92, 8'd99, 8'd138, 8'd129, 8'd96, 8'd136, 8'd77, 8'd101, 8'd69, 8'd65, 8'd156, 8'd119, 8'd166, 8'd176, 8'd167, 8'd130, 8'd161, 8'd69, 8'd142, 8'd69, 8'd130, 8'd65, 8'd88, 8'd128, 8'd78, 8'd84, 8'd137, 8'd88, 8'd129, 8'd81, 8'd109, 8'd146, 8'd94, 8'd153, 8'd167, 8'd124, 8'd155, 8'd80, 8'd119, 8'd80, 8'd62, 8'd134, 8'd99, 8'd129, 8'd73, 8'd120, 8'd83, 8'd85, 8'd137, 8'd106, 8'd134, 8'd119, 8'd109, 8'd137, 8'd120, 8'd134, 8'd68, 8'd109, 8'd127, 8'd100, 8'd156, 8'd103, 8'd157, 8'd80, 8'd143, 8'd131, 8'd157, 8'd90, 8'd149, 8'd85, 8'd133, 8'd134, 8'd74, 8'd161, 8'd143, 8'd125, 8'd160, 8'd109, 8'd81, 8'd154, 8'd100, 8'd96, 8'd114, 8'd124, 8'd95, 8'd107, 8'd43, 8'd81, 8'd77, 8'd120, 8'd129, 8'd137, 8'd143, 8'd98, 8'd107, 8'd90, 8'd125, 8'd99, 8'd76, 8'd143, 8'd64, 8'd98, 8'd139, 8'd136, 8'd134, 8'd85, 8'd83, 8'd105, 8'd145, 8'd87, 8'd87, 8'd70, 8'd112, 8'd79, 8'd106, 8'd120, 8'd85, 8'd147, 8'd109, 8'd75, 8'd61, 8'd63, 8'd65, 8'd113, 8'd116, 8'd106, 8'd66, 8'd132, 8'd83, 8'd147, 8'd84, 8'd109, 8'd143, 8'd96, 8'd85, 8'd148, 8'd65, 8'd116, 8'd123, 8'd108, 8'd88, 8'd76, 8'd90, 8'd157, 8'd137, 8'd139, 8'd96, 8'd139, 8'd129, 8'd149, 8'd161, 8'd120, 8'd148, 8'd135, 8'd108, 8'd76, 8'd137, 8'd89, 8'd89, 8'd145, 8'd139, 8'd182, 8'd125, 8'd114, 8'd92, 8'd117, 8'd82, 8'd132, 8'd77, 8'd112, 8'd53, 8'd122, 8'd102, 8'd93, 8'd120, 8'd117, 8'd92, 8'd89, 8'd96, 8'd126, 8'd104, 8'd105, 8'd160, 8'd111, 8'd99, 8'd72, 8'd107, 8'd137, 8'd73, 8'd159, 8'd129, 8'd145, 8'd121, 8'd161, 8'd62, 8'd66, 8'd76, 8'd72, 8'd92, 8'd137, 8'd153, 8'd140, 8'd92, 8'd72, 8'd122, 8'd136, 8'd127, 8'd152, 8'd143, 8'd91, 8'd133, 8'd164, 8'd87, 8'd118, 8'd136, 8'd96, 8'd82, 8'd160, 8'd86, 8'd114, 8'd90, 8'd118, 8'd142, 8'd132, 8'd121, 8'd110, 8'd94, 8'd134, 8'd108, 8'd103, 8'd92, 8'd83, 8'd59, 8'd57, 8'd118, 8'd120, 8'd110, 8'd119, 8'd68, 8'd152, 8'd82, 8'd88, 8'd158, 8'd120, 8'd107, 8'd100, 8'd154, 8'd94, 8'd101, 8'd87, 8'd67, 8'd106, 8'd138, 8'd147, 8'd64, 8'd150, 8'd121, 8'd158, 8'd110, 8'd41, 8'd52, 8'd122, 8'd143, 8'd167, 8'd104, 8'd151, 8'd146, 8'd158, 8'd133, 8'd130, 8'd145, 8'd146, 8'd71, 8'd157, 8'd114, 8'd111, 8'd116, 8'd117, 8'd80, 8'd71, 8'd71, 8'd109, 8'd130, 8'd131, 8'd138, 8'd100, 8'd73, 8'd49, 8'd90, 8'd99, 8'd91, 8'd136, 8'd152, 8'd88, 8'd125, 8'd75, 8'd70, 8'd129, 8'd79, 8'd108, 8'd86, 8'd111, 8'd74, 8'd68, 8'd83, 8'd81, 8'd156, 8'd157, 8'd92, 8'd142, 8'd137, 8'd164, 8'd132, 8'd101, 8'd78, 8'd89, 8'd136, 8'd123, 8'd135, 8'd100, 8'd152, 8'd134, 8'd168, 8'd156, 8'd148, 8'd117, 8'd167, 8'd96, 8'd101, 8'd63, 8'd158, 8'd149, 8'd114, 8'd163, 8'd93, 8'd145, 8'd147, 8'd136, 8'd89, 8'd94, 8'd133, 8'd163, 8'd135, 8'd51, 8'd74, 8'd75, 8'd177, 8'd171, 8'd110, 8'd144, 8'd90, 8'd122, 8'd113, 8'd72, 8'd157, 8'd152, 8'd93, 8'd114, 8'd101, 8'd113, 8'd177, 8'd159, 8'd125, 8'd188, 8'd181, 8'd190, 8'd180, 8'd127, 8'd130, 8'd142, 8'd144, 8'd143, 8'd137, 8'd180, 8'd117, 8'd153, 8'd119, 8'd163, 8'd152, 8'd137, 8'd114, 8'd131, 8'd97, 8'd176, 8'd111, 8'd143, 8'd149, 8'd145, 8'd161, 8'd159, 8'd130, 8'd176, 8'd97, 8'd105, 8'd73, 8'd135, 8'd177, 8'd116, 8'd142, 8'd154, 8'd148, 8'd116, 8'd145, 8'd83, 8'd135, 8'd82, 8'd121, 8'd118, 8'd53, 8'd93, 8'd80, 8'd126, 8'd185, 8'd122, 8'd182, 8'd131, 8'd93, 8'd132, 8'd120, 8'd151, 8'd69, 8'd109, 8'd144, 8'd77, 8'd106, 8'd151, 8'd177, 8'd117, 8'd98, 8'd156, 8'd89, 8'd133, 8'd146, 8'd55, 8'd99, 8'd108, 8'd145, 8'd86, 8'd143, 8'd175, 8'd98, 8'd116, 8'd112, 8'd96, 8'd84, 8'd81, 8'd127, 8'd110, 8'd71, 8'd136, 8'd102, 8'd77, 8'd179, 8'd141, 8'd122, 8'd86, 8'd85, 8'd117, 8'd112, 8'd155, 8'd117, 8'd99, 8'd147, 8'd69, 8'd120, 8'd165, 8'd121, 8'd140, 8'd85, 8'd94, 8'd145, 8'd92, 8'd143, 8'd143, 8'd95, 8'd70, 8'd83, 8'd47, 8'd86, 8'd77, 8'd149, 8'd88, 8'd134, 8'd112, 8'd87, 8'd153, 8'd94, 8'd150, 8'd134, 8'd135, 8'd100, 8'd161, 8'd161, 8'd107, 8'd114, 8'd159, 8'd172, 8'd123, 8'd120, 8'd109, 8'd110, 8'd86, 8'd156, 8'd137, 8'd83, 8'd70, 8'd58, 8'd90, 8'd65, 8'd109, 8'd131, 8'd69, 8'd105, 8'd80, 8'd97, 8'd154, 8'd109, 8'd81, 8'd112, 8'd89, 8'd158, 8'd122, 8'd95, 8'd147, 8'd128, 8'd178, 8'd167, 8'd153, 8'd149, 8'd118, 8'd76, 8'd52, 8'd104, 8'd54, 8'd65, 8'd83, 8'd102, 8'd147, 8'd100, 8'd149, 8'd86, 8'd100, 8'd172, 8'd164, 8'd141, 8'd143, 8'd117, 8'd140, 8'd130, 8'd108, 8'd125, 8'd107, 8'd144, 8'd168, 8'd153, 8'd115, 8'd123, 8'd80, 8'd143, 8'd104, 8'd75, 8'd106, 8'd95, 8'd93, 8'd111, 8'd114, 8'd172, 8'd139, 8'd164, 8'd107, 8'd116, 8'd136, 8'd119, 8'd149, 8'd94, 8'd135, 8'd121, 8'd99, 8'd88, 8'd142, 8'd88, 8'd132, 8'd144, 8'd92, 8'd77, 8'd85, 8'd115, 8'd83, 8'd119, 8'd141, 8'd109, 8'd149, 8'd159, 8'd114, 8'd103, 8'd120, 8'd77, 8'd118, 8'd161, 8'd147, 8'd140, 8'd187, 8'd106, 8'd176, 8'd117, 8'd129, 8'd82, 8'd123, 8'd85, 8'd58, 8'd160, 8'd93, 8'd156, 8'd98, 8'd121, 8'd118, 8'd142, 8'd136, 8'd117, 8'd130, 8'd145, 8'd133, 8'd103, 8'd91, 8'd106, 8'd152, 8'd188, 8'd158, 8'd105, 8'd187, 8'd166, 8'd173, 8'd137, 8'd134, 8'd172, 8'd150, 8'd138, 8'd136, 8'd154, 8'd188, 8'd153, 8'd95, 8'd167, 8'd152, 8'd91, 8'd154, 8'd103, 8'd173, 8'd99, 8'd144, 8'd126, 8'd149, 8'd97, 8'd95, 8'd124, 8'd164, 8'd142, 8'd113, 8'd139, 8'd184, 8'd93, 8'd67, 8'd137, 8'd109, 8'd133, 8'd161, 8'd164, 8'd101, 8'd167, 8'd122, 8'd173, 8'd179, 8'd169, 8'd109, 8'd120, 8'd112, 8'd167, 8'd130, 8'd146, 8'd120, 8'd132, 8'd90, 8'd138, 8'd140, 8'd105, 8'd73, 8'd136, 8'd82, 8'd158, 8'd107, 8'd126, 8'd131, 8'd169, 8'd142, 8'd85, 8'd132, 8'd131, 8'd151, 8'd166, 8'd80, 8'd139, 8'd124, 8'd90, 8'd150, 8'd93, 8'd81})
) cell_0_14 (
    .clk(clk),
    .input_index(index_0_13_14),
    .input_value(value_0_13_14),
    .input_result(result_0_13_14),
    .input_enable(enable_0_13_14),
    .output_index(index_0_14_15),
    .output_value(value_0_14_15),
    .output_result(result_0_14_15),
    .output_enable(enable_0_14_15)
);

wire [10-1:0] index_0_15_16;
wire [`DATA_WIDTH-1:0] value_0_15_16;
wire [`DATA_WIDTH*4:0] result_0_15_16;
wire enable_0_15_16;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd159, 8'd170, 8'd87, 8'd99, 8'd154, 8'd123, 8'd171, 8'd172, 8'd98, 8'd125, 8'd119, 8'd102, 8'd165, 8'd191, 8'd164, 8'd89, 8'd89, 8'd173, 8'd137, 8'd164, 8'd156, 8'd124, 8'd81, 8'd131, 8'd155, 8'd162, 8'd99, 8'd165, 8'd141, 8'd70, 8'd108, 8'd82, 8'd173, 8'd102, 8'd151, 8'd151, 8'd172, 8'd150, 8'd172, 8'd149, 8'd178, 8'd180, 8'd146, 8'd164, 8'd174, 8'd187, 8'd186, 8'd113, 8'd130, 8'd168, 8'd177, 8'd177, 8'd99, 8'd84, 8'd136, 8'd167, 8'd116, 8'd95, 8'd156, 8'd129, 8'd87, 8'd151, 8'd172, 8'd131, 8'd180, 8'd98, 8'd132, 8'd175, 8'd182, 8'd121, 8'd178, 8'd94, 8'd124, 8'd107, 8'd162, 8'd123, 8'd113, 8'd101, 8'd74, 8'd119, 8'd79, 8'd85, 8'd114, 8'd163, 8'd127, 8'd131, 8'd78, 8'd101, 8'd101, 8'd111, 8'd133, 8'd184, 8'd99, 8'd131, 8'd141, 8'd95, 8'd84, 8'd159, 8'd85, 8'd106, 8'd159, 8'd105, 8'd129, 8'd134, 8'd149, 8'd78, 8'd95, 8'd51, 8'd122, 8'd153, 8'd74, 8'd125, 8'd125, 8'd62, 8'd134, 8'd97, 8'd181, 8'd110, 8'd165, 8'd149, 8'd104, 8'd144, 8'd74, 8'd124, 8'd120, 8'd105, 8'd91, 8'd119, 8'd80, 8'd128, 8'd98, 8'd128, 8'd78, 8'd131, 8'd163, 8'd76, 8'd48, 8'd90, 8'd96, 8'd129, 8'd107, 8'd68, 8'd97, 8'd147, 8'd164, 8'd85, 8'd108, 8'd101, 8'd74, 8'd82, 8'd80, 8'd92, 8'd146, 8'd125, 8'd131, 8'd118, 8'd143, 8'd89, 8'd128, 8'd108, 8'd116, 8'd102, 8'd142, 8'd72, 8'd141, 8'd123, 8'd103, 8'd147, 8'd123, 8'd127, 8'd165, 8'd144, 8'd128, 8'd132, 8'd81, 8'd151, 8'd132, 8'd94, 8'd106, 8'd91, 8'd137, 8'd68, 8'd82, 8'd162, 8'd147, 8'd94, 8'd176, 8'd129, 8'd104, 8'd177, 8'd157, 8'd74, 8'd85, 8'd151, 8'd109, 8'd76, 8'd118, 8'd98, 8'd110, 8'd102, 8'd160, 8'd122, 8'd81, 8'd127, 8'd116, 8'd86, 8'd128, 8'd133, 8'd113, 8'd112, 8'd72, 8'd95, 8'd155, 8'd131, 8'd127, 8'd158, 8'd176, 8'd173, 8'd116, 8'd66, 8'd61, 8'd129, 8'd167, 8'd112, 8'd85, 8'd124, 8'd135, 8'd183, 8'd157, 8'd120, 8'd136, 8'd87, 8'd108, 8'd117, 8'd90, 8'd112, 8'd154, 8'd130, 8'd168, 8'd111, 8'd84, 8'd120, 8'd159, 8'd103, 8'd161, 8'd161, 8'd109, 8'd113, 8'd75, 8'd147, 8'd125, 8'd141, 8'd137, 8'd133, 8'd103, 8'd85, 8'd135, 8'd84, 8'd82, 8'd112, 8'd72, 8'd147, 8'd111, 8'd107, 8'd70, 8'd169, 8'd103, 8'd125, 8'd84, 8'd163, 8'd138, 8'd70, 8'd142, 8'd78, 8'd146, 8'd83, 8'd76, 8'd87, 8'd142, 8'd166, 8'd182, 8'd97, 8'd174, 8'd138, 8'd161, 8'd127, 8'd124, 8'd121, 8'd82, 8'd59, 8'd129, 8'd113, 8'd79, 8'd129, 8'd118, 8'd115, 8'd76, 8'd133, 8'd79, 8'd62, 8'd145, 8'd96, 8'd97, 8'd183, 8'd137, 8'd104, 8'd128, 8'd119, 8'd135, 8'd180, 8'd140, 8'd152, 8'd118, 8'd149, 8'd101, 8'd102, 8'd128, 8'd130, 8'd126, 8'd141, 8'd147, 8'd163, 8'd149, 8'd113, 8'd78, 8'd93, 8'd110, 8'd113, 8'd140, 8'd110, 8'd125, 8'd161, 8'd80, 8'd83, 8'd116, 8'd158, 8'd126, 8'd184, 8'd116, 8'd82, 8'd70, 8'd106, 8'd107, 8'd75, 8'd140, 8'd158, 8'd64, 8'd59, 8'd80, 8'd95, 8'd100, 8'd96, 8'd94, 8'd61, 8'd144, 8'd65, 8'd123, 8'd98, 8'd75, 8'd132, 8'd118, 8'd86, 8'd130, 8'd139, 8'd103, 8'd140, 8'd93, 8'd90, 8'd40, 8'd86, 8'd148, 8'd72, 8'd71, 8'd141, 8'd120, 8'd132, 8'd85, 8'd114, 8'd82, 8'd114, 8'd52, 8'd119, 8'd92, 8'd65, 8'd64, 8'd128, 8'd111, 8'd160, 8'd156, 8'd99, 8'd109, 8'd145, 8'd124, 8'd114, 8'd157, 8'd119, 8'd69, 8'd118, 8'd106, 8'd98, 8'd147, 8'd144, 8'd71, 8'd92, 8'd155, 8'd140, 8'd60, 8'd24, 8'd96, 8'd51, 8'd84, 8'd93, 8'd69, 8'd103, 8'd110, 8'd109, 8'd115, 8'd171, 8'd93, 8'd146, 8'd114, 8'd110, 8'd73, 8'd81, 8'd142, 8'd127, 8'd168, 8'd101, 8'd129, 8'd139, 8'd167, 8'd73, 8'd95, 8'd180, 8'd62, 8'd100, 8'd67, 8'd67, 8'd138, 8'd83, 8'd63, 8'd103, 8'd176, 8'd138, 8'd182, 8'd107, 8'd161, 8'd165, 8'd75, 8'd161, 8'd125, 8'd94, 8'd143, 8'd105, 8'd172, 8'd128, 8'd110, 8'd135, 8'd166, 8'd122, 8'd129, 8'd131, 8'd149, 8'd135, 8'd102, 8'd81, 8'd101, 8'd98, 8'd140, 8'd101, 8'd122, 8'd158, 8'd132, 8'd122, 8'd168, 8'd165, 8'd75, 8'd128, 8'd63, 8'd53, 8'd163, 8'd163, 8'd105, 8'd111, 8'd84, 8'd159, 8'd104, 8'd159, 8'd208, 8'd109, 8'd122, 8'd135, 8'd124, 8'd154, 8'd145, 8'd165, 8'd151, 8'd98, 8'd166, 8'd176, 8'd157, 8'd115, 8'd140, 8'd136, 8'd174, 8'd155, 8'd80, 8'd103, 8'd151, 8'd138, 8'd156, 8'd101, 8'd87, 8'd99, 8'd181, 8'd116, 8'd196, 8'd193, 8'd120, 8'd130, 8'd150, 8'd104, 8'd155, 8'd164, 8'd170, 8'd143, 8'd89, 8'd121, 8'd160, 8'd134, 8'd117, 8'd146, 8'd142, 8'd159, 8'd138, 8'd101, 8'd125, 8'd146, 8'd143, 8'd135, 8'd176, 8'd141, 8'd155, 8'd170, 8'd204, 8'd166, 8'd173, 8'd98, 8'd111, 8'd136, 8'd102, 8'd146, 8'd83, 8'd148, 8'd85, 8'd143, 8'd93, 8'd156, 8'd110, 8'd125, 8'd112, 8'd94, 8'd73, 8'd121, 8'd75, 8'd144, 8'd145, 8'd153, 8'd167, 8'd177, 8'd118, 8'd198, 8'd165, 8'd122, 8'd161, 8'd139, 8'd146, 8'd105, 8'd105, 8'd107, 8'd93, 8'd155, 8'd111, 8'd100, 8'd131, 8'd110, 8'd115, 8'd142, 8'd80, 8'd104, 8'd149, 8'd85, 8'd84, 8'd118, 8'd119, 8'd166, 8'd100, 8'd162, 8'd106, 8'd113, 8'd151, 8'd115, 8'd96, 8'd120, 8'd115, 8'd145, 8'd109, 8'd134, 8'd58, 8'd132, 8'd139, 8'd87, 8'd84, 8'd156, 8'd161, 8'd138, 8'd118, 8'd131, 8'd144, 8'd77, 8'd79, 8'd93, 8'd117, 8'd131, 8'd118, 8'd55, 8'd64, 8'd91, 8'd128, 8'd139, 8'd105, 8'd87, 8'd98, 8'd70, 8'd67, 8'd139, 8'd141, 8'd66, 8'd129, 8'd63, 8'd66, 8'd105, 8'd152, 8'd99, 8'd98, 8'd115, 8'd98, 8'd116, 8'd92, 8'd132, 8'd89, 8'd74, 8'd107, 8'd148, 8'd132, 8'd94, 8'd154, 8'd120, 8'd166, 8'd141, 8'd78, 8'd80, 8'd93, 8'd133, 8'd145, 8'd131, 8'd118, 8'd71, 8'd77, 8'd86, 8'd154, 8'd110, 8'd115, 8'd135, 8'd98, 8'd77, 8'd117, 8'd48, 8'd53, 8'd67, 8'd82, 8'd77, 8'd105, 8'd80, 8'd132, 8'd113, 8'd111, 8'd76, 8'd101, 8'd69, 8'd95, 8'd134, 8'd66, 8'd151, 8'd124, 8'd133, 8'd86, 8'd165, 8'd126, 8'd109, 8'd102, 8'd82, 8'd87, 8'd75, 8'd81, 8'd136, 8'd110, 8'd59, 8'd72, 8'd113, 8'd86, 8'd134, 8'd156, 8'd117, 8'd99, 8'd110, 8'd113, 8'd70, 8'd79, 8'd141, 8'd119, 8'd112, 8'd65, 8'd132, 8'd126, 8'd131, 8'd88, 8'd96, 8'd76, 8'd105, 8'd119, 8'd159, 8'd175, 8'd171, 8'd103, 8'd125, 8'd144, 8'd74, 8'd143, 8'd121, 8'd154, 8'd119, 8'd154, 8'd124, 8'd167, 8'd83, 8'd114, 8'd84, 8'd142, 8'd154, 8'd150, 8'd116, 8'd165, 8'd115, 8'd140, 8'd113, 8'd115, 8'd116, 8'd143, 8'd166, 8'd98, 8'd141, 8'd80, 8'd162, 8'd92, 8'd128, 8'd73, 8'd127, 8'd119, 8'd86, 8'd125, 8'd143, 8'd97, 8'd93, 8'd169, 8'd105, 8'd154, 8'd72, 8'd162, 8'd168, 8'd158, 8'd170, 8'd132, 8'd135})
) cell_0_15 (
    .clk(clk),
    .input_index(index_0_14_15),
    .input_value(value_0_14_15),
    .input_result(result_0_14_15),
    .input_enable(enable_0_14_15),
    .output_index(index_0_15_16),
    .output_value(value_0_15_16),
    .output_result(result_0_15_16),
    .output_enable(enable_0_15_16)
);

wire [10-1:0] index_0_16_17;
wire [`DATA_WIDTH-1:0] value_0_16_17;
wire [`DATA_WIDTH*4:0] result_0_16_17;
wire enable_0_16_17;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd109, 8'd107, 8'd155, 8'd156, 8'd105, 8'd154, 8'd102, 8'd85, 8'd156, 8'd115, 8'd132, 8'd173, 8'd142, 8'd210, 8'd197, 8'd103, 8'd118, 8'd187, 8'd92, 8'd94, 8'd176, 8'd98, 8'd80, 8'd98, 8'd101, 8'd88, 8'd108, 8'd127, 8'd139, 8'd155, 8'd153, 8'd97, 8'd98, 8'd184, 8'd166, 8'd153, 8'd129, 8'd185, 8'd136, 8'd176, 8'd180, 8'd130, 8'd165, 8'd133, 8'd179, 8'd209, 8'd188, 8'd171, 8'd171, 8'd144, 8'd118, 8'd90, 8'd73, 8'd84, 8'd169, 8'd148, 8'd95, 8'd158, 8'd156, 8'd74, 8'd152, 8'd116, 8'd162, 8'd162, 8'd195, 8'd204, 8'd142, 8'd192, 8'd158, 8'd188, 8'd181, 8'd149, 8'd167, 8'd120, 8'd194, 8'd163, 8'd175, 8'd156, 8'd110, 8'd109, 8'd76, 8'd149, 8'd158, 8'd140, 8'd137, 8'd67, 8'd128, 8'd62, 8'd113, 8'd151, 8'd143, 8'd133, 8'd143, 8'd151, 8'd151, 8'd116, 8'd82, 8'd159, 8'd137, 8'd89, 8'd90, 8'd113, 8'd113, 8'd119, 8'd94, 8'd189, 8'd176, 8'd144, 8'd144, 8'd122, 8'd155, 8'd72, 8'd143, 8'd109, 8'd90, 8'd131, 8'd74, 8'd96, 8'd104, 8'd120, 8'd88, 8'd182, 8'd144, 8'd148, 8'd175, 8'd116, 8'd69, 8'd65, 8'd112, 8'd105, 8'd158, 8'd152, 8'd120, 8'd104, 8'd104, 8'd148, 8'd138, 8'd128, 8'd82, 8'd142, 8'd96, 8'd111, 8'd159, 8'd151, 8'd59, 8'd144, 8'd128, 8'd103, 8'd94, 8'd110, 8'd96, 8'd100, 8'd72, 8'd112, 8'd51, 8'd149, 8'd130, 8'd90, 8'd131, 8'd96, 8'd172, 8'd160, 8'd152, 8'd161, 8'd141, 8'd109, 8'd134, 8'd132, 8'd84, 8'd137, 8'd137, 8'd146, 8'd76, 8'd121, 8'd95, 8'd89, 8'd128, 8'd114, 8'd109, 8'd127, 8'd66, 8'd124, 8'd61, 8'd54, 8'd76, 8'd137, 8'd75, 8'd153, 8'd96, 8'd101, 8'd69, 8'd122, 8'd139, 8'd102, 8'd158, 8'd150, 8'd110, 8'd83, 8'd104, 8'd152, 8'd140, 8'd122, 8'd146, 8'd93, 8'd121, 8'd138, 8'd139, 8'd113, 8'd127, 8'd162, 8'd89, 8'd79, 8'd65, 8'd93, 8'd106, 8'd87, 8'd119, 8'd65, 8'd126, 8'd116, 8'd106, 8'd120, 8'd105, 8'd74, 8'd128, 8'd93, 8'd94, 8'd110, 8'd72, 8'd62, 8'd123, 8'd93, 8'd157, 8'd106, 8'd95, 8'd145, 8'd65, 8'd92, 8'd94, 8'd71, 8'd143, 8'd74, 8'd51, 8'd134, 8'd71, 8'd79, 8'd80, 8'd73, 8'd175, 8'd126, 8'd144, 8'd148, 8'd180, 8'd149, 8'd80, 8'd72, 8'd59, 8'd84, 8'd160, 8'd134, 8'd90, 8'd76, 8'd127, 8'd106, 8'd153, 8'd112, 8'd117, 8'd115, 8'd154, 8'd119, 8'd121, 8'd53, 8'd54, 8'd103, 8'd115, 8'd130, 8'd131, 8'd119, 8'd127, 8'd103, 8'd113, 8'd103, 8'd69, 8'd133, 8'd136, 8'd65, 8'd129, 8'd125, 8'd138, 8'd88, 8'd127, 8'd75, 8'd125, 8'd164, 8'd165, 8'd83, 8'd149, 8'd74, 8'd118, 8'd86, 8'd122, 8'd72, 8'd65, 8'd137, 8'd174, 8'd153, 8'd175, 8'd112, 8'd152, 8'd158, 8'd84, 8'd76, 8'd80, 8'd70, 8'd156, 8'd134, 8'd153, 8'd110, 8'd110, 8'd152, 8'd158, 8'd179, 8'd140, 8'd113, 8'd59, 8'd54, 8'd35, 8'd92, 8'd49, 8'd66, 8'd86, 8'd146, 8'd126, 8'd163, 8'd172, 8'd170, 8'd89, 8'd161, 8'd155, 8'd41, 8'd102, 8'd74, 8'd151, 8'd132, 8'd110, 8'd122, 8'd136, 8'd126, 8'd166, 8'd160, 8'd105, 8'd64, 8'd49, 8'd75, 8'd22, 8'd48, 8'd116, 8'd66, 8'd74, 8'd152, 8'd144, 8'd96, 8'd81, 8'd157, 8'd134, 8'd165, 8'd114, 8'd41, 8'd65, 8'd50, 8'd68, 8'd76, 8'd83, 8'd168, 8'd132, 8'd200, 8'd151, 8'd119, 8'd175, 8'd135, 8'd104, 8'd62, 8'd51, 8'd58, 8'd73, 8'd106, 8'd131, 8'd101, 8'd120, 8'd169, 8'd133, 8'd83, 8'd159, 8'd145, 8'd94, 8'd134, 8'd114, 8'd93, 8'd68, 8'd112, 8'd123, 8'd151, 8'd134, 8'd141, 8'd123, 8'd170, 8'd145, 8'd121, 8'd81, 8'd86, 8'd63, 8'd92, 8'd94, 8'd114, 8'd87, 8'd119, 8'd131, 8'd95, 8'd142, 8'd145, 8'd138, 8'd95, 8'd123, 8'd118, 8'd90, 8'd160, 8'd165, 8'd138, 8'd167, 8'd102, 8'd137, 8'd177, 8'd208, 8'd149, 8'd103, 8'd104, 8'd127, 8'd49, 8'd146, 8'd104, 8'd91, 8'd100, 8'd186, 8'd155, 8'd206, 8'd148, 8'd153, 8'd129, 8'd80, 8'd73, 8'd95, 8'd93, 8'd108, 8'd134, 8'd88, 8'd156, 8'd129, 8'd116, 8'd152, 8'd176, 8'd138, 8'd211, 8'd153, 8'd137, 8'd97, 8'd121, 8'd133, 8'd95, 8'd94, 8'd82, 8'd95, 8'd197, 8'd139, 8'd186, 8'd142, 8'd156, 8'd116, 8'd132, 8'd123, 8'd18, 8'd88, 8'd92, 8'd93, 8'd158, 8'd184, 8'd116, 8'd180, 8'd121, 8'd154, 8'd152, 8'd147, 8'd120, 8'd109, 8'd164, 8'd167, 8'd103, 8'd158, 8'd96, 8'd115, 8'd191, 8'd160, 8'd122, 8'd177, 8'd160, 8'd97, 8'd119, 8'd52, 8'd116, 8'd41, 8'd108, 8'd70, 8'd138, 8'd100, 8'd141, 8'd100, 8'd94, 8'd106, 8'd188, 8'd155, 8'd102, 8'd114, 8'd119, 8'd160, 8'd97, 8'd126, 8'd122, 8'd101, 8'd139, 8'd146, 8'd111, 8'd169, 8'd148, 8'd143, 8'd155, 8'd86, 8'd48, 8'd132, 8'd82, 8'd136, 8'd141, 8'd107, 8'd116, 8'd132, 8'd121, 8'd190, 8'd162, 8'd130, 8'd95, 8'd164, 8'd178, 8'd141, 8'd164, 8'd127, 8'd116, 8'd154, 8'd195, 8'd154, 8'd172, 8'd85, 8'd110, 8'd105, 8'd146, 8'd145, 8'd108, 8'd131, 8'd101, 8'd77, 8'd97, 8'd147, 8'd81, 8'd165, 8'd167, 8'd146, 8'd179, 8'd140, 8'd182, 8'd161, 8'd95, 8'd128, 8'd128, 8'd145, 8'd109, 8'd140, 8'd135, 8'd167, 8'd133, 8'd152, 8'd85, 8'd110, 8'd112, 8'd79, 8'd119, 8'd84, 8'd78, 8'd139, 8'd124, 8'd83, 8'd151, 8'd133, 8'd148, 8'd90, 8'd107, 8'd151, 8'd125, 8'd126, 8'd125, 8'd111, 8'd99, 8'd126, 8'd132, 8'd127, 8'd123, 8'd144, 8'd100, 8'd119, 8'd142, 8'd144, 8'd77, 8'd133, 8'd61, 8'd57, 8'd92, 8'd99, 8'd122, 8'd139, 8'd137, 8'd92, 8'd115, 8'd123, 8'd94, 8'd105, 8'd153, 8'd134, 8'd107, 8'd135, 8'd123, 8'd164, 8'd130, 8'd108, 8'd113, 8'd91, 8'd172, 8'd118, 8'd99, 8'd71, 8'd104, 8'd77, 8'd99, 8'd80, 8'd97, 8'd119, 8'd101, 8'd156, 8'd126, 8'd131, 8'd149, 8'd162, 8'd166, 8'd155, 8'd138, 8'd110, 8'd74, 8'd154, 8'd131, 8'd131, 8'd137, 8'd114, 8'd154, 8'd162, 8'd149, 8'd107, 8'd96, 8'd128, 8'd158, 8'd77, 8'd129, 8'd151, 8'd56, 8'd131, 8'd125, 8'd100, 8'd96, 8'd154, 8'd149, 8'd95, 8'd64, 8'd120, 8'd124, 8'd95, 8'd132, 8'd108, 8'd108, 8'd155, 8'd96, 8'd174, 8'd150, 8'd111, 8'd147, 8'd73, 8'd145, 8'd142, 8'd116, 8'd163, 8'd138, 8'd76, 8'd122, 8'd64, 8'd109, 8'd143, 8'd147, 8'd108, 8'd182, 8'd114, 8'd179, 8'd80, 8'd110, 8'd152, 8'd129, 8'd131, 8'd64, 8'd82, 8'd96, 8'd162, 8'd74, 8'd107, 8'd116, 8'd88, 8'd157, 8'd113, 8'd152, 8'd154, 8'd85, 8'd140, 8'd168, 8'd114, 8'd84, 8'd94, 8'd140, 8'd107, 8'd119, 8'd166, 8'd128, 8'd96, 8'd111, 8'd71, 8'd86, 8'd132, 8'd113, 8'd177, 8'd104, 8'd69, 8'd107, 8'd154, 8'd169, 8'd151, 8'd128, 8'd88, 8'd162, 8'd102, 8'd81, 8'd102, 8'd90, 8'd77, 8'd132, 8'd90, 8'd93, 8'd130, 8'd74, 8'd78, 8'd85, 8'd116, 8'd113, 8'd103, 8'd134, 8'd137, 8'd122, 8'd105, 8'd105, 8'd144, 8'd72, 8'd146, 8'd78, 8'd71, 8'd101})
) cell_0_16 (
    .clk(clk),
    .input_index(index_0_15_16),
    .input_value(value_0_15_16),
    .input_result(result_0_15_16),
    .input_enable(enable_0_15_16),
    .output_index(index_0_16_17),
    .output_value(value_0_16_17),
    .output_result(result_0_16_17),
    .output_enable(enable_0_16_17)
);

wire [10-1:0] index_0_17_18;
wire [`DATA_WIDTH-1:0] value_0_17_18;
wire [`DATA_WIDTH*4:0] result_0_17_18;
wire enable_0_17_18;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd88, 8'd104, 8'd114, 8'd132, 8'd123, 8'd126, 8'd93, 8'd85, 8'd47, 8'd68, 8'd100, 8'd56, 8'd127, 8'd137, 8'd114, 8'd124, 8'd55, 8'd53, 8'd95, 8'd122, 8'd142, 8'd60, 8'd67, 8'd156, 8'd130, 8'd124, 8'd104, 8'd132, 8'd85, 8'd149, 8'd78, 8'd78, 8'd161, 8'd152, 8'd97, 8'd73, 8'd34, 8'd49, 8'd124, 8'd89, 8'd117, 8'd131, 8'd53, 8'd93, 8'd128, 8'd79, 8'd71, 8'd140, 8'd150, 8'd155, 8'd130, 8'd158, 8'd99, 8'd78, 8'd86, 8'd143, 8'd137, 8'd163, 8'd102, 8'd144, 8'd111, 8'd68, 8'd142, 8'd82, 8'd81, 8'd91, 8'd91, 8'd119, 8'd83, 8'd167, 8'd149, 8'd72, 8'd94, 8'd142, 8'd163, 8'd94, 8'd169, 8'd105, 8'd137, 8'd120, 8'd99, 8'd147, 8'd141, 8'd89, 8'd98, 8'd90, 8'd90, 8'd150, 8'd137, 8'd152, 8'd181, 8'd133, 8'd126, 8'd128, 8'd98, 8'd162, 8'd99, 8'd111, 8'd79, 8'd165, 8'd146, 8'd173, 8'd95, 8'd133, 8'd126, 8'd151, 8'd125, 8'd157, 8'd81, 8'd97, 8'd97, 8'd110, 8'd130, 8'd176, 8'd95, 8'd132, 8'd167, 8'd158, 8'd178, 8'd144, 8'd122, 8'd155, 8'd179, 8'd113, 8'd77, 8'd143, 8'd104, 8'd108, 8'd116, 8'd137, 8'd168, 8'd142, 8'd92, 8'd114, 8'd117, 8'd130, 8'd122, 8'd83, 8'd148, 8'd82, 8'd115, 8'd164, 8'd138, 8'd119, 8'd178, 8'd109, 8'd154, 8'd167, 8'd115, 8'd135, 8'd151, 8'd94, 8'd131, 8'd64, 8'd100, 8'd126, 8'd132, 8'd107, 8'd108, 8'd138, 8'd157, 8'd109, 8'd110, 8'd108, 8'd157, 8'd169, 8'd103, 8'd173, 8'd154, 8'd84, 8'd116, 8'd125, 8'd122, 8'd163, 8'd142, 8'd131, 8'd151, 8'd122, 8'd110, 8'd107, 8'd120, 8'd77, 8'd62, 8'd44, 8'd78, 8'd127, 8'd131, 8'd73, 8'd150, 8'd136, 8'd73, 8'd92, 8'd99, 8'd103, 8'd94, 8'd119, 8'd101, 8'd138, 8'd103, 8'd169, 8'd76, 8'd137, 8'd163, 8'd102, 8'd88, 8'd141, 8'd114, 8'd80, 8'd110, 8'd105, 8'd48, 8'd40, 8'd63, 8'd104, 8'd122, 8'd144, 8'd126, 8'd141, 8'd86, 8'd127, 8'd161, 8'd92, 8'd83, 8'd124, 8'd177, 8'd105, 8'd131, 8'd144, 8'd109, 8'd152, 8'd103, 8'd96, 8'd153, 8'd64, 8'd115, 8'd137, 8'd135, 8'd149, 8'd112, 8'd120, 8'd63, 8'd56, 8'd123, 8'd72, 8'd112, 8'd118, 8'd94, 8'd170, 8'd162, 8'd111, 8'd88, 8'd113, 8'd88, 8'd116, 8'd146, 8'd150, 8'd129, 8'd58, 8'd69, 8'd143, 8'd73, 8'd118, 8'd90, 8'd109, 8'd85, 8'd149, 8'd143, 8'd68, 8'd78, 8'd123, 8'd64, 8'd67, 8'd103, 8'd110, 8'd127, 8'd130, 8'd146, 8'd157, 8'd132, 8'd127, 8'd73, 8'd174, 8'd76, 8'd122, 8'd141, 8'd60, 8'd68, 8'd99, 8'd166, 8'd169, 8'd121, 8'd174, 8'd129, 8'd119, 8'd123, 8'd122, 8'd105, 8'd75, 8'd58, 8'd132, 8'd112, 8'd80, 8'd113, 8'd96, 8'd77, 8'd89, 8'd90, 8'd133, 8'd147, 8'd138, 8'd150, 8'd106, 8'd73, 8'd113, 8'd79, 8'd80, 8'd80, 8'd160, 8'd132, 8'd160, 8'd190, 8'd141, 8'd179, 8'd108, 8'd92, 8'd65, 8'd98, 8'd129, 8'd98, 8'd144, 8'd140, 8'd144, 8'd94, 8'd109, 8'd135, 8'd122, 8'd107, 8'd117, 8'd112, 8'd138, 8'd94, 8'd79, 8'd89, 8'd110, 8'd151, 8'd94, 8'd185, 8'd118, 8'd124, 8'd160, 8'd134, 8'd164, 8'd80, 8'd99, 8'd139, 8'd100, 8'd141, 8'd132, 8'd164, 8'd160, 8'd152, 8'd105, 8'd91, 8'd164, 8'd91, 8'd140, 8'd91, 8'd135, 8'd83, 8'd65, 8'd96, 8'd84, 8'd179, 8'd165, 8'd118, 8'd169, 8'd98, 8'd169, 8'd105, 8'd97, 8'd84, 8'd145, 8'd119, 8'd106, 8'd76, 8'd96, 8'd150, 8'd119, 8'd105, 8'd139, 8'd125, 8'd154, 8'd127, 8'd134, 8'd158, 8'd110, 8'd47, 8'd145, 8'd95, 8'd87, 8'd183, 8'd159, 8'd129, 8'd188, 8'd113, 8'd143, 8'd137, 8'd163, 8'd163, 8'd94, 8'd156, 8'd159, 8'd170, 8'd113, 8'd127, 8'd142, 8'd86, 8'd97, 8'd151, 8'd123, 8'd88, 8'd100, 8'd122, 8'd72, 8'd96, 8'd89, 8'd144, 8'd125, 8'd135, 8'd161, 8'd130, 8'd118, 8'd140, 8'd149, 8'd87, 8'd170, 8'd174, 8'd177, 8'd110, 8'd88, 8'd84, 8'd153, 8'd146, 8'd148, 8'd107, 8'd134, 8'd108, 8'd130, 8'd123, 8'd129, 8'd155, 8'd94, 8'd104, 8'd117, 8'd98, 8'd115, 8'd163, 8'd182, 8'd184, 8'd162, 8'd190, 8'd125, 8'd109, 8'd125, 8'd127, 8'd126, 8'd95, 8'd85, 8'd110, 8'd78, 8'd148, 8'd82, 8'd146, 8'd88, 8'd147, 8'd149, 8'd107, 8'd170, 8'd167, 8'd97, 8'd126, 8'd120, 8'd100, 8'd122, 8'd167, 8'd124, 8'd101, 8'd124, 8'd158, 8'd113, 8'd69, 8'd156, 8'd157, 8'd86, 8'd90, 8'd82, 8'd148, 8'd134, 8'd150, 8'd151, 8'd101, 8'd132, 8'd128, 8'd104, 8'd127, 8'd155, 8'd173, 8'd125, 8'd61, 8'd131, 8'd83, 8'd174, 8'd165, 8'd87, 8'd120, 8'd123, 8'd167, 8'd84, 8'd77, 8'd104, 8'd72, 8'd122, 8'd150, 8'd108, 8'd166, 8'd133, 8'd124, 8'd140, 8'd102, 8'd93, 8'd73, 8'd130, 8'd134, 8'd107, 8'd153, 8'd113, 8'd150, 8'd122, 8'd124, 8'd169, 8'd96, 8'd93, 8'd135, 8'd105, 8'd67, 8'd99, 8'd76, 8'd100, 8'd118, 8'd151, 8'd163, 8'd80, 8'd112, 8'd154, 8'd147, 8'd144, 8'd119, 8'd67, 8'd81, 8'd122, 8'd162, 8'd97, 8'd109, 8'd76, 8'd105, 8'd100, 8'd123, 8'd79, 8'd92, 8'd136, 8'd165, 8'd127, 8'd155, 8'd104, 8'd103, 8'd102, 8'd90, 8'd142, 8'd99, 8'd151, 8'd80, 8'd101, 8'd157, 8'd182, 8'd142, 8'd137, 8'd101, 8'd154, 8'd118, 8'd180, 8'd143, 8'd119, 8'd154, 8'd81, 8'd146, 8'd125, 8'd144, 8'd85, 8'd145, 8'd154, 8'd114, 8'd125, 8'd125, 8'd108, 8'd143, 8'd159, 8'd130, 8'd144, 8'd92, 8'd108, 8'd149, 8'd110, 8'd161, 8'd97, 8'd120, 8'd102, 8'd82, 8'd81, 8'd120, 8'd112, 8'd151, 8'd115, 8'd96, 8'd87, 8'd70, 8'd79, 8'd84, 8'd111, 8'd161, 8'd110, 8'd140, 8'd156, 8'd93, 8'd101, 8'd170, 8'd94, 8'd162, 8'd151, 8'd165, 8'd174, 8'd91, 8'd169, 8'd120, 8'd117, 8'd136, 8'd111, 8'd138, 8'd121, 8'd134, 8'd125, 8'd62, 8'd107, 8'd103, 8'd87, 8'd95, 8'd86, 8'd63, 8'd93, 8'd131, 8'd96, 8'd142, 8'd159, 8'd120, 8'd111, 8'd151, 8'd159, 8'd165, 8'd101, 8'd151, 8'd148, 8'd74, 8'd117, 8'd109, 8'd160, 8'd103, 8'd126, 8'd48, 8'd87, 8'd113, 8'd83, 8'd115, 8'd46, 8'd79, 8'd116, 8'd100, 8'd79, 8'd89, 8'd71, 8'd79, 8'd61, 8'd137, 8'd102, 8'd76, 8'd64, 8'd82, 8'd96, 8'd161, 8'd78, 8'd121, 8'd87, 8'd142, 8'd117, 8'd88, 8'd79, 8'd131, 8'd124, 8'd131, 8'd108, 8'd61, 8'd114, 8'd69, 8'd138, 8'd87, 8'd73, 8'd41, 8'd101, 8'd103, 8'd66, 8'd59, 8'd134, 8'd122, 8'd84, 8'd119, 8'd91, 8'd88, 8'd141, 8'd130, 8'd125, 8'd106, 8'd151, 8'd154, 8'd94, 8'd146, 8'd66, 8'd98, 8'd68, 8'd148, 8'd59, 8'd118, 8'd71, 8'd102, 8'd106, 8'd64, 8'd47, 8'd128, 8'd92, 8'd139, 8'd82, 8'd96, 8'd80, 8'd115, 8'd97, 8'd145, 8'd76, 8'd114, 8'd131, 8'd103, 8'd164, 8'd91, 8'd142, 8'd108, 8'd169, 8'd138, 8'd159, 8'd102, 8'd131, 8'd158, 8'd162, 8'd121, 8'd153, 8'd132, 8'd80, 8'd80, 8'd132, 8'd122, 8'd101, 8'd132, 8'd80, 8'd146, 8'd147, 8'd78, 8'd146, 8'd139, 8'd156})
) cell_0_17 (
    .clk(clk),
    .input_index(index_0_16_17),
    .input_value(value_0_16_17),
    .input_result(result_0_16_17),
    .input_enable(enable_0_16_17),
    .output_index(index_0_17_18),
    .output_value(value_0_17_18),
    .output_result(result_0_17_18),
    .output_enable(enable_0_17_18)
);

wire [10-1:0] index_0_18_19;
wire [`DATA_WIDTH-1:0] value_0_18_19;
wire [`DATA_WIDTH*4:0] result_0_18_19;
wire enable_0_18_19;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd94, 8'd170, 8'd167, 8'd116, 8'd162, 8'd142, 8'd147, 8'd122, 8'd126, 8'd127, 8'd162, 8'd124, 8'd93, 8'd76, 8'd181, 8'd111, 8'd138, 8'd114, 8'd142, 8'd95, 8'd130, 8'd133, 8'd177, 8'd149, 8'd110, 8'd168, 8'd142, 8'd114, 8'd96, 8'd96, 8'd172, 8'd134, 8'd164, 8'd107, 8'd125, 8'd99, 8'd67, 8'd121, 8'd84, 8'd71, 8'd123, 8'd130, 8'd111, 8'd108, 8'd144, 8'd77, 8'd126, 8'd127, 8'd77, 8'd89, 8'd117, 8'd57, 8'd102, 8'd168, 8'd93, 8'd102, 8'd110, 8'd77, 8'd136, 8'd86, 8'd91, 8'd138, 8'd88, 8'd99, 8'd60, 8'd93, 8'd101, 8'd113, 8'd119, 8'd146, 8'd83, 8'd156, 8'd149, 8'd121, 8'd111, 8'd125, 8'd160, 8'd80, 8'd140, 8'd139, 8'd102, 8'd88, 8'd100, 8'd130, 8'd168, 8'd138, 8'd149, 8'd112, 8'd94, 8'd125, 8'd135, 8'd156, 8'd90, 8'd142, 8'd105, 8'd126, 8'd133, 8'd103, 8'd138, 8'd141, 8'd114, 8'd109, 8'd160, 8'd162, 8'd159, 8'd179, 8'd112, 8'd95, 8'd164, 8'd172, 8'd93, 8'd114, 8'd145, 8'd92, 8'd140, 8'd105, 8'd56, 8'd134, 8'd133, 8'd164, 8'd108, 8'd91, 8'd151, 8'd151, 8'd88, 8'd166, 8'd139, 8'd131, 8'd133, 8'd131, 8'd104, 8'd129, 8'd136, 8'd97, 8'd144, 8'd114, 8'd187, 8'd87, 8'd96, 8'd71, 8'd105, 8'd147, 8'd142, 8'd121, 8'd132, 8'd66, 8'd125, 8'd85, 8'd98, 8'd171, 8'd144, 8'd166, 8'd126, 8'd153, 8'd152, 8'd85, 8'd81, 8'd115, 8'd141, 8'd77, 8'd122, 8'd123, 8'd85, 8'd180, 8'd175, 8'd176, 8'd89, 8'd141, 8'd159, 8'd117, 8'd129, 8'd55, 8'd91, 8'd149, 8'd143, 8'd81, 8'd160, 8'd112, 8'd103, 8'd156, 8'd165, 8'd159, 8'd162, 8'd143, 8'd146, 8'd145, 8'd147, 8'd155, 8'd147, 8'd127, 8'd148, 8'd124, 8'd107, 8'd170, 8'd98, 8'd88, 8'd175, 8'd132, 8'd106, 8'd84, 8'd131, 8'd101, 8'd133, 8'd109, 8'd73, 8'd132, 8'd104, 8'd156, 8'd96, 8'd120, 8'd76, 8'd111, 8'd127, 8'd124, 8'd123, 8'd129, 8'd168, 8'd126, 8'd118, 8'd158, 8'd150, 8'd155, 8'd144, 8'd76, 8'd154, 8'd142, 8'd48, 8'd95, 8'd75, 8'd161, 8'd134, 8'd77, 8'd168, 8'd109, 8'd172, 8'd127, 8'd164, 8'd97, 8'd135, 8'd100, 8'd136, 8'd111, 8'd153, 8'd123, 8'd154, 8'd80, 8'd119, 8'd88, 8'd169, 8'd140, 8'd77, 8'd84, 8'd129, 8'd155, 8'd76, 8'd102, 8'd155, 8'd103, 8'd99, 8'd164, 8'd172, 8'd145, 8'd73, 8'd81, 8'd160, 8'd84, 8'd100, 8'd86, 8'd125, 8'd64, 8'd135, 8'd145, 8'd72, 8'd167, 8'd150, 8'd125, 8'd179, 8'd145, 8'd157, 8'd68, 8'd109, 8'd101, 8'd87, 8'd116, 8'd141, 8'd95, 8'd134, 8'd75, 8'd86, 8'd173, 8'd142, 8'd121, 8'd92, 8'd101, 8'd160, 8'd96, 8'd98, 8'd45, 8'd95, 8'd80, 8'd128, 8'd70, 8'd157, 8'd84, 8'd125, 8'd101, 8'd120, 8'd111, 8'd101, 8'd95, 8'd106, 8'd69, 8'd110, 8'd142, 8'd84, 8'd166, 8'd87, 8'd159, 8'd72, 8'd71, 8'd97, 8'd104, 8'd174, 8'd165, 8'd65, 8'd108, 8'd60, 8'd124, 8'd135, 8'd69, 8'd91, 8'd84, 8'd104, 8'd182, 8'd149, 8'd166, 8'd127, 8'd54, 8'd77, 8'd145, 8'd161, 8'd160, 8'd76, 8'd83, 8'd116, 8'd88, 8'd159, 8'd159, 8'd154, 8'd138, 8'd151, 8'd116, 8'd87, 8'd77, 8'd111, 8'd135, 8'd90, 8'd72, 8'd95, 8'd130, 8'd91, 8'd146, 8'd163, 8'd88, 8'd108, 8'd128, 8'd63, 8'd82, 8'd124, 8'd158, 8'd157, 8'd80, 8'd76, 8'd143, 8'd133, 8'd84, 8'd179, 8'd184, 8'd119, 8'd105, 8'd111, 8'd78, 8'd165, 8'd160, 8'd68, 8'd66, 8'd121, 8'd156, 8'd159, 8'd178, 8'd150, 8'd175, 8'd122, 8'd108, 8'd134, 8'd149, 8'd103, 8'd56, 8'd85, 8'd143, 8'd149, 8'd128, 8'd87, 8'd169, 8'd106, 8'd175, 8'd180, 8'd172, 8'd163, 8'd87, 8'd135, 8'd104, 8'd95, 8'd128, 8'd120, 8'd152, 8'd106, 8'd120, 8'd115, 8'd99, 8'd94, 8'd96, 8'd135, 8'd127, 8'd61, 8'd59, 8'd123, 8'd94, 8'd96, 8'd108, 8'd101, 8'd148, 8'd186, 8'd104, 8'd112, 8'd165, 8'd177, 8'd107, 8'd78, 8'd155, 8'd83, 8'd92, 8'd128, 8'd148, 8'd175, 8'd92, 8'd145, 8'd101, 8'd135, 8'd120, 8'd175, 8'd119, 8'd69, 8'd61, 8'd121, 8'd119, 8'd126, 8'd97, 8'd83, 8'd105, 8'd137, 8'd157, 8'd189, 8'd138, 8'd170, 8'd130, 8'd131, 8'd133, 8'd75, 8'd148, 8'd113, 8'd167, 8'd188, 8'd98, 8'd121, 8'd155, 8'd155, 8'd196, 8'd160, 8'd183, 8'd128, 8'd148, 8'd127, 8'd100, 8'd155, 8'd137, 8'd126, 8'd108, 8'd160, 8'd90, 8'd135, 8'd97, 8'd86, 8'd149, 8'd122, 8'd99, 8'd85, 8'd103, 8'd77, 8'd170, 8'd147, 8'd149, 8'd161, 8'd98, 8'd89, 8'd177, 8'd137, 8'd175, 8'd150, 8'd96, 8'd179, 8'd109, 8'd85, 8'd130, 8'd136, 8'd156, 8'd143, 8'd65, 8'd74, 8'd121, 8'd96, 8'd116, 8'd125, 8'd96, 8'd114, 8'd167, 8'd124, 8'd135, 8'd155, 8'd111, 8'd157, 8'd85, 8'd113, 8'd100, 8'd167, 8'd121, 8'd85, 8'd146, 8'd97, 8'd102, 8'd138, 8'd103, 8'd99, 8'd65, 8'd126, 8'd72, 8'd112, 8'd86, 8'd154, 8'd105, 8'd122, 8'd139, 8'd154, 8'd140, 8'd165, 8'd135, 8'd181, 8'd84, 8'd132, 8'd78, 8'd175, 8'd144, 8'd209, 8'd116, 8'd94, 8'd133, 8'd103, 8'd124, 8'd126, 8'd129, 8'd72, 8'd87, 8'd53, 8'd50, 8'd76, 8'd103, 8'd130, 8'd85, 8'd136, 8'd156, 8'd111, 8'd130, 8'd190, 8'd142, 8'd155, 8'd65, 8'd181, 8'd167, 8'd153, 8'd198, 8'd185, 8'd109, 8'd184, 8'd104, 8'd120, 8'd157, 8'd102, 8'd131, 8'd69, 8'd71, 8'd85, 8'd111, 8'd137, 8'd132, 8'd104, 8'd83, 8'd129, 8'd113, 8'd109, 8'd148, 8'd91, 8'd98, 8'd150, 8'd161, 8'd129, 8'd93, 8'd111, 8'd137, 8'd127, 8'd191, 8'd120, 8'd127, 8'd162, 8'd96, 8'd125, 8'd169, 8'd90, 8'd147, 8'd83, 8'd133, 8'd69, 8'd145, 8'd77, 8'd102, 8'd166, 8'd96, 8'd125, 8'd112, 8'd153, 8'd175, 8'd121, 8'd143, 8'd80, 8'd132, 8'd65, 8'd166, 8'd120, 8'd153, 8'd146, 8'd166, 8'd91, 8'd159, 8'd165, 8'd167, 8'd168, 8'd80, 8'd115, 8'd145, 8'd113, 8'd178, 8'd140, 8'd140, 8'd163, 8'd108, 8'd120, 8'd154, 8'd103, 8'd97, 8'd88, 8'd145, 8'd94, 8'd107, 8'd125, 8'd81, 8'd69, 8'd138, 8'd98, 8'd85, 8'd152, 8'd172, 8'd79, 8'd115, 8'd161, 8'd90, 8'd121, 8'd128, 8'd120, 8'd116, 8'd132, 8'd98, 8'd72, 8'd93, 8'd130, 8'd165, 8'd163, 8'd97, 8'd131, 8'd103, 8'd107, 8'd152, 8'd81, 8'd104, 8'd117, 8'd73, 8'd103, 8'd144, 8'd60, 8'd104, 8'd121, 8'd97, 8'd150, 8'd102, 8'd80, 8'd122, 8'd119, 8'd123, 8'd88, 8'd47, 8'd58, 8'd102, 8'd142, 8'd108, 8'd108, 8'd147, 8'd68, 8'd73, 8'd168, 8'd88, 8'd119, 8'd122, 8'd117, 8'd170, 8'd72, 8'd136, 8'd102, 8'd115, 8'd92, 8'd125, 8'd94, 8'd146, 8'd137, 8'd85, 8'd58, 8'd137, 8'd149, 8'd82, 8'd102, 8'd81, 8'd121, 8'd88, 8'd106, 8'd153, 8'd114, 8'd101, 8'd170, 8'd158, 8'd82, 8'd147, 8'd127, 8'd166, 8'd123, 8'd80, 8'd156, 8'd104, 8'd127, 8'd151, 8'd124, 8'd130, 8'd117, 8'd74, 8'd155, 8'd145, 8'd150, 8'd85, 8'd88, 8'd152, 8'd116, 8'd98, 8'd131, 8'd145, 8'd115, 8'd164, 8'd76, 8'd74})
) cell_0_18 (
    .clk(clk),
    .input_index(index_0_17_18),
    .input_value(value_0_17_18),
    .input_result(result_0_17_18),
    .input_enable(enable_0_17_18),
    .output_index(index_0_18_19),
    .output_value(value_0_18_19),
    .output_result(result_0_18_19),
    .output_enable(enable_0_18_19)
);

wire [10-1:0] index_0_19_20;
wire [`DATA_WIDTH-1:0] value_0_19_20;
wire [`DATA_WIDTH*4:0] result_0_19_20;
wire enable_0_19_20;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd100, 8'd70, 8'd86, 8'd90, 8'd127, 8'd136, 8'd141, 8'd98, 8'd93, 8'd97, 8'd152, 8'd160, 8'd190, 8'd122, 8'd108, 8'd157, 8'd140, 8'd137, 8'd82, 8'd119, 8'd126, 8'd91, 8'd85, 8'd107, 8'd104, 8'd98, 8'd96, 8'd92, 8'd141, 8'd106, 8'd77, 8'd100, 8'd78, 8'd152, 8'd166, 8'd77, 8'd97, 8'd106, 8'd150, 8'd123, 8'd145, 8'd82, 8'd134, 8'd78, 8'd88, 8'd163, 8'd94, 8'd144, 8'd142, 8'd73, 8'd129, 8'd80, 8'd109, 8'd137, 8'd99, 8'd105, 8'd153, 8'd163, 8'd149, 8'd91, 8'd139, 8'd105, 8'd146, 8'd113, 8'd145, 8'd68, 8'd140, 8'd126, 8'd135, 8'd92, 8'd112, 8'd128, 8'd156, 8'd164, 8'd165, 8'd127, 8'd139, 8'd122, 8'd154, 8'd123, 8'd98, 8'd95, 8'd129, 8'd141, 8'd161, 8'd87, 8'd153, 8'd104, 8'd75, 8'd124, 8'd63, 8'd119, 8'd67, 8'd97, 8'd128, 8'd134, 8'd137, 8'd129, 8'd90, 8'd142, 8'd152, 8'd135, 8'd100, 8'd78, 8'd98, 8'd153, 8'd125, 8'd145, 8'd169, 8'd83, 8'd133, 8'd92, 8'd139, 8'd106, 8'd158, 8'd101, 8'd118, 8'd66, 8'd55, 8'd148, 8'd128, 8'd124, 8'd90, 8'd86, 8'd150, 8'd144, 8'd108, 8'd124, 8'd91, 8'd138, 8'd159, 8'd123, 8'd185, 8'd161, 8'd165, 8'd156, 8'd77, 8'd139, 8'd117, 8'd83, 8'd109, 8'd134, 8'd55, 8'd61, 8'd50, 8'd88, 8'd79, 8'd75, 8'd72, 8'd117, 8'd160, 8'd156, 8'd112, 8'd79, 8'd134, 8'd97, 8'd116, 8'd66, 8'd135, 8'd97, 8'd152, 8'd91, 8'd169, 8'd146, 8'd99, 8'd75, 8'd137, 8'd90, 8'd122, 8'd151, 8'd84, 8'd86, 8'd93, 8'd27, 8'd132, 8'd70, 8'd72, 8'd132, 8'd69, 8'd69, 8'd130, 8'd143, 8'd97, 8'd90, 8'd126, 8'd117, 8'd75, 8'd109, 8'd133, 8'd77, 8'd57, 8'd125, 8'd121, 8'd102, 8'd113, 8'd144, 8'd127, 8'd121, 8'd134, 8'd56, 8'd75, 8'd106, 8'd39, 8'd128, 8'd73, 8'd78, 8'd122, 8'd106, 8'd131, 8'd102, 8'd124, 8'd139, 8'd109, 8'd112, 8'd115, 8'd40, 8'd55, 8'd78, 8'd47, 8'd109, 8'd158, 8'd71, 8'd144, 8'd169, 8'd128, 8'd74, 8'd113, 8'd75, 8'd99, 8'd100, 8'd101, 8'd133, 8'd110, 8'd92, 8'd51, 8'd145, 8'd132, 8'd119, 8'd105, 8'd123, 8'd51, 8'd78, 8'd121, 8'd63, 8'd114, 8'd121, 8'd120, 8'd128, 8'd134, 8'd92, 8'd150, 8'd97, 8'd115, 8'd171, 8'd63, 8'd117, 8'd36, 8'd88, 8'd115, 8'd110, 8'd140, 8'd83, 8'd50, 8'd137, 8'd136, 8'd155, 8'd110, 8'd73, 8'd81, 8'd96, 8'd136, 8'd46, 8'd100, 8'd133, 8'd102, 8'd88, 8'd83, 8'd121, 8'd145, 8'd133, 8'd71, 8'd85, 8'd92, 8'd46, 8'd91, 8'd54, 8'd140, 8'd110, 8'd151, 8'd161, 8'd110, 8'd105, 8'd142, 8'd170, 8'd107, 8'd77, 8'd78, 8'd52, 8'd150, 8'd104, 8'd88, 8'd92, 8'd128, 8'd151, 8'd79, 8'd147, 8'd102, 8'd100, 8'd103, 8'd89, 8'd88, 8'd111, 8'd80, 8'd151, 8'd85, 8'd148, 8'd165, 8'd166, 8'd159, 8'd127, 8'd87, 8'd165, 8'd158, 8'd121, 8'd85, 8'd134, 8'd124, 8'd153, 8'd180, 8'd129, 8'd131, 8'd125, 8'd65, 8'd171, 8'd119, 8'd90, 8'd116, 8'd122, 8'd37, 8'd117, 8'd165, 8'd110, 8'd133, 8'd172, 8'd144, 8'd140, 8'd93, 8'd82, 8'd107, 8'd134, 8'd109, 8'd80, 8'd89, 8'd133, 8'd124, 8'd137, 8'd139, 8'd163, 8'd148, 8'd120, 8'd163, 8'd170, 8'd93, 8'd139, 8'd73, 8'd132, 8'd103, 8'd77, 8'd131, 8'd179, 8'd86, 8'd148, 8'd167, 8'd118, 8'd129, 8'd106, 8'd76, 8'd133, 8'd126, 8'd69, 8'd45, 8'd98, 8'd145, 8'd104, 8'd101, 8'd170, 8'd134, 8'd145, 8'd156, 8'd152, 8'd128, 8'd71, 8'd96, 8'd141, 8'd100, 8'd59, 8'd94, 8'd157, 8'd105, 8'd166, 8'd114, 8'd162, 8'd93, 8'd129, 8'd123, 8'd142, 8'd46, 8'd78, 8'd112, 8'd160, 8'd164, 8'd189, 8'd172, 8'd112, 8'd96, 8'd175, 8'd97, 8'd194, 8'd112, 8'd85, 8'd83, 8'd128, 8'd51, 8'd82, 8'd104, 8'd154, 8'd155, 8'd108, 8'd159, 8'd162, 8'd140, 8'd137, 8'd116, 8'd131, 8'd68, 8'd69, 8'd125, 8'd124, 8'd168, 8'd117, 8'd127, 8'd141, 8'd119, 8'd164, 8'd125, 8'd148, 8'd119, 8'd93, 8'd154, 8'd30, 8'd82, 8'd9, 8'd117, 8'd112, 8'd169, 8'd169, 8'd104, 8'd140, 8'd156, 8'd112, 8'd188, 8'd167, 8'd119, 8'd74, 8'd75, 8'd93, 8'd165, 8'd85, 8'd137, 8'd138, 8'd107, 8'd146, 8'd145, 8'd147, 8'd107, 8'd164, 8'd110, 8'd117, 8'd80, 8'd30, 8'd90, 8'd136, 8'd89, 8'd83, 8'd105, 8'd148, 8'd126, 8'd162, 8'd211, 8'd113, 8'd174, 8'd99, 8'd99, 8'd66, 8'd127, 8'd124, 8'd121, 8'd150, 8'd111, 8'd136, 8'd97, 8'd166, 8'd88, 8'd143, 8'd162, 8'd119, 8'd108, 8'd27, 8'd95, 8'd126, 8'd151, 8'd86, 8'd173, 8'd128, 8'd141, 8'd122, 8'd171, 8'd124, 8'd128, 8'd133, 8'd92, 8'd134, 8'd107, 8'd77, 8'd82, 8'd101, 8'd134, 8'd88, 8'd170, 8'd127, 8'd186, 8'd98, 8'd100, 8'd87, 8'd63, 8'd83, 8'd74, 8'd115, 8'd93, 8'd94, 8'd82, 8'd161, 8'd157, 8'd170, 8'd87, 8'd117, 8'd122, 8'd131, 8'd79, 8'd140, 8'd127, 8'd119, 8'd144, 8'd135, 8'd166, 8'd150, 8'd194, 8'd175, 8'd167, 8'd104, 8'd78, 8'd67, 8'd37, 8'd60, 8'd87, 8'd112, 8'd148, 8'd97, 8'd164, 8'd152, 8'd130, 8'd71, 8'd51, 8'd128, 8'd148, 8'd75, 8'd135, 8'd87, 8'd137, 8'd100, 8'd151, 8'd81, 8'd124, 8'd159, 8'd118, 8'd153, 8'd102, 8'd79, 8'd99, 8'd90, 8'd131, 8'd81, 8'd147, 8'd116, 8'd82, 8'd97, 8'd125, 8'd97, 8'd112, 8'd116, 8'd38, 8'd67, 8'd104, 8'd91, 8'd65, 8'd142, 8'd99, 8'd156, 8'd152, 8'd181, 8'd151, 8'd121, 8'd129, 8'd138, 8'd168, 8'd74, 8'd164, 8'd142, 8'd87, 8'd90, 8'd126, 8'd176, 8'd89, 8'd113, 8'd130, 8'd149, 8'd72, 8'd59, 8'd45, 8'd94, 8'd107, 8'd100, 8'd113, 8'd79, 8'd72, 8'd92, 8'd169, 8'd147, 8'd132, 8'd185, 8'd161, 8'd139, 8'd123, 8'd123, 8'd105, 8'd153, 8'd155, 8'd92, 8'd97, 8'd111, 8'd183, 8'd174, 8'd132, 8'd73, 8'd138, 8'd130, 8'd110, 8'd59, 8'd100, 8'd107, 8'd54, 8'd27, 8'd130, 8'd119, 8'd102, 8'd137, 8'd142, 8'd148, 8'd155, 8'd108, 8'd82, 8'd102, 8'd161, 8'd90, 8'd84, 8'd75, 8'd106, 8'd99, 8'd72, 8'd117, 8'd147, 8'd79, 8'd135, 8'd83, 8'd73, 8'd43, 8'd16, 8'd6, 8'd84, 8'd62, 8'd76, 8'd92, 8'd61, 8'd110, 8'd107, 8'd62, 8'd128, 8'd109, 8'd153, 8'd75, 8'd154, 8'd142, 8'd153, 8'd150, 8'd68, 8'd76, 8'd98, 8'd118, 8'd51, 8'd125, 8'd67, 8'd125, 8'd130, 8'd140, 8'd133, 8'd109, 8'd101, 8'd23, 8'd25, 8'd71, 8'd100, 8'd62, 8'd129, 8'd75, 8'd105, 8'd78, 8'd139, 8'd127, 8'd167, 8'd162, 8'd141, 8'd91, 8'd77, 8'd60, 8'd88, 8'd147, 8'd103, 8'd80, 8'd50, 8'd138, 8'd104, 8'd117, 8'd53, 8'd53, 8'd75, 8'd91, 8'd140, 8'd153, 8'd85, 8'd68, 8'd87, 8'd96, 8'd152, 8'd134, 8'd83, 8'd114, 8'd126, 8'd80, 8'd131, 8'd103, 8'd135, 8'd141, 8'd144, 8'd118, 8'd119, 8'd122, 8'd72, 8'd76, 8'd71, 8'd107, 8'd73, 8'd155, 8'd134, 8'd146, 8'd132, 8'd99, 8'd97, 8'd151, 8'd141, 8'd155, 8'd92, 8'd107, 8'd91, 8'd150})
) cell_0_19 (
    .clk(clk),
    .input_index(index_0_18_19),
    .input_value(value_0_18_19),
    .input_result(result_0_18_19),
    .input_enable(enable_0_18_19),
    .output_index(index_0_19_20),
    .output_value(value_0_19_20),
    .output_result(result_0_19_20),
    .output_enable(enable_0_19_20)
);

wire [10-1:0] index_0_20_21;
wire [`DATA_WIDTH-1:0] value_0_20_21;
wire [`DATA_WIDTH*4:0] result_0_20_21;
wire enable_0_20_21;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd86, 8'd84, 8'd85, 8'd110, 8'd89, 8'd147, 8'd105, 8'd116, 8'd59, 8'd92, 8'd83, 8'd102, 8'd89, 8'd107, 8'd146, 8'd110, 8'd112, 8'd155, 8'd111, 8'd139, 8'd58, 8'd76, 8'd77, 8'd92, 8'd125, 8'd99, 8'd165, 8'd170, 8'd100, 8'd70, 8'd97, 8'd164, 8'd121, 8'd114, 8'd157, 8'd91, 8'd161, 8'd139, 8'd145, 8'd121, 8'd169, 8'd146, 8'd155, 8'd154, 8'd99, 8'd182, 8'd117, 8'd82, 8'd92, 8'd134, 8'd170, 8'd167, 8'd127, 8'd116, 8'd144, 8'd114, 8'd149, 8'd71, 8'd165, 8'd102, 8'd175, 8'd141, 8'd180, 8'd109, 8'd85, 8'd141, 8'd162, 8'd95, 8'd120, 8'd133, 8'd103, 8'd99, 8'd114, 8'd86, 8'd140, 8'd94, 8'd97, 8'd161, 8'd111, 8'd168, 8'd79, 8'd86, 8'd90, 8'd133, 8'd86, 8'd151, 8'd86, 8'd99, 8'd181, 8'd187, 8'd179, 8'd141, 8'd71, 8'd134, 8'd124, 8'd100, 8'd75, 8'd151, 8'd142, 8'd145, 8'd86, 8'd86, 8'd129, 8'd117, 8'd141, 8'd158, 8'd136, 8'd111, 8'd67, 8'd161, 8'd110, 8'd143, 8'd93, 8'd71, 8'd107, 8'd98, 8'd123, 8'd115, 8'd171, 8'd110, 8'd154, 8'd59, 8'd131, 8'd114, 8'd156, 8'd120, 8'd79, 8'd128, 8'd107, 8'd166, 8'd151, 8'd156, 8'd149, 8'd147, 8'd82, 8'd103, 8'd75, 8'd114, 8'd101, 8'd73, 8'd158, 8'd119, 8'd139, 8'd149, 8'd182, 8'd154, 8'd145, 8'd146, 8'd60, 8'd84, 8'd108, 8'd106, 8'd131, 8'd146, 8'd84, 8'd141, 8'd128, 8'd123, 8'd139, 8'd72, 8'd67, 8'd66, 8'd107, 8'd75, 8'd68, 8'd121, 8'd166, 8'd120, 8'd170, 8'd164, 8'd157, 8'd121, 8'd146, 8'd99, 8'd77, 8'd121, 8'd86, 8'd94, 8'd82, 8'd98, 8'd91, 8'd112, 8'd72, 8'd130, 8'd74, 8'd104, 8'd88, 8'd76, 8'd74, 8'd57, 8'd103, 8'd165, 8'd118, 8'd80, 8'd82, 8'd119, 8'd144, 8'd95, 8'd111, 8'd109, 8'd113, 8'd103, 8'd88, 8'd97, 8'd118, 8'd82, 8'd117, 8'd122, 8'd75, 8'd154, 8'd128, 8'd87, 8'd144, 8'd126, 8'd132, 8'd137, 8'd104, 8'd154, 8'd80, 8'd152, 8'd138, 8'd90, 8'd147, 8'd157, 8'd157, 8'd71, 8'd168, 8'd121, 8'd157, 8'd106, 8'd71, 8'd149, 8'd112, 8'd99, 8'd131, 8'd76, 8'd132, 8'd91, 8'd146, 8'd143, 8'd95, 8'd89, 8'd137, 8'd79, 8'd96, 8'd132, 8'd127, 8'd69, 8'd73, 8'd153, 8'd148, 8'd120, 8'd140, 8'd128, 8'd154, 8'd131, 8'd71, 8'd127, 8'd107, 8'd84, 8'd124, 8'd80, 8'd113, 8'd87, 8'd171, 8'd163, 8'd105, 8'd164, 8'd75, 8'd97, 8'd129, 8'd78, 8'd81, 8'd154, 8'd109, 8'd99, 8'd79, 8'd131, 8'd78, 8'd155, 8'd68, 8'd98, 8'd95, 8'd159, 8'd68, 8'd138, 8'd140, 8'd131, 8'd89, 8'd118, 8'd158, 8'd145, 8'd162, 8'd110, 8'd104, 8'd132, 8'd110, 8'd137, 8'd154, 8'd155, 8'd84, 8'd143, 8'd140, 8'd80, 8'd64, 8'd142, 8'd148, 8'd140, 8'd93, 8'd164, 8'd131, 8'd79, 8'd157, 8'd104, 8'd156, 8'd131, 8'd154, 8'd155, 8'd174, 8'd174, 8'd129, 8'd60, 8'd65, 8'd138, 8'd111, 8'd145, 8'd125, 8'd192, 8'd91, 8'd143, 8'd163, 8'd79, 8'd123, 8'd143, 8'd109, 8'd127, 8'd147, 8'd73, 8'd114, 8'd76, 8'd101, 8'd91, 8'd115, 8'd83, 8'd139, 8'd142, 8'd136, 8'd166, 8'd109, 8'd100, 8'd103, 8'd83, 8'd143, 8'd122, 8'd197, 8'd156, 8'd138, 8'd180, 8'd123, 8'd156, 8'd119, 8'd120, 8'd88, 8'd109, 8'd89, 8'd74, 8'd120, 8'd114, 8'd146, 8'd107, 8'd97, 8'd112, 8'd144, 8'd106, 8'd140, 8'd150, 8'd65, 8'd96, 8'd136, 8'd157, 8'd99, 8'd137, 8'd138, 8'd192, 8'd178, 8'd151, 8'd158, 8'd196, 8'd150, 8'd77, 8'd127, 8'd127, 8'd85, 8'd93, 8'd122, 8'd103, 8'd106, 8'd126, 8'd150, 8'd162, 8'd179, 8'd139, 8'd145, 8'd137, 8'd115, 8'd119, 8'd118, 8'd152, 8'd105, 8'd178, 8'd116, 8'd99, 8'd166, 8'd118, 8'd174, 8'd99, 8'd88, 8'd122, 8'd111, 8'd136, 8'd90, 8'd124, 8'd102, 8'd75, 8'd79, 8'd143, 8'd152, 8'd146, 8'd119, 8'd73, 8'd117, 8'd66, 8'd127, 8'd87, 8'd107, 8'd119, 8'd154, 8'd186, 8'd108, 8'd115, 8'd185, 8'd159, 8'd90, 8'd83, 8'd91, 8'd115, 8'd123, 8'd141, 8'd89, 8'd107, 8'd90, 8'd113, 8'd127, 8'd117, 8'd75, 8'd149, 8'd95, 8'd87, 8'd129, 8'd104, 8'd151, 8'd134, 8'd115, 8'd173, 8'd160, 8'd182, 8'd180, 8'd138, 8'd178, 8'd108, 8'd128, 8'd126, 8'd103, 8'd130, 8'd65, 8'd124, 8'd99, 8'd154, 8'd155, 8'd138, 8'd158, 8'd156, 8'd149, 8'd117, 8'd89, 8'd149, 8'd123, 8'd85, 8'd139, 8'd146, 8'd160, 8'd186, 8'd160, 8'd157, 8'd151, 8'd114, 8'd107, 8'd152, 8'd131, 8'd39, 8'd99, 8'd138, 8'd108, 8'd153, 8'd151, 8'd137, 8'd112, 8'd139, 8'd129, 8'd169, 8'd80, 8'd113, 8'd148, 8'd81, 8'd82, 8'd122, 8'd88, 8'd72, 8'd93, 8'd175, 8'd155, 8'd161, 8'd139, 8'd127, 8'd62, 8'd146, 8'd76, 8'd64, 8'd105, 8'd67, 8'd159, 8'd85, 8'd147, 8'd80, 8'd152, 8'd171, 8'd178, 8'd169, 8'd109, 8'd76, 8'd78, 8'd125, 8'd87, 8'd92, 8'd116, 8'd97, 8'd79, 8'd68, 8'd121, 8'd153, 8'd164, 8'd123, 8'd76, 8'd135, 8'd118, 8'd65, 8'd105, 8'd70, 8'd113, 8'd156, 8'd135, 8'd107, 8'd156, 8'd94, 8'd178, 8'd90, 8'd149, 8'd74, 8'd120, 8'd110, 8'd164, 8'd77, 8'd156, 8'd161, 8'd89, 8'd138, 8'd100, 8'd84, 8'd97, 8'd96, 8'd144, 8'd112, 8'd118, 8'd54, 8'd86, 8'd99, 8'd98, 8'd150, 8'd161, 8'd95, 8'd98, 8'd113, 8'd146, 8'd133, 8'd103, 8'd165, 8'd105, 8'd155, 8'd110, 8'd131, 8'd93, 8'd127, 8'd141, 8'd165, 8'd82, 8'd157, 8'd105, 8'd96, 8'd139, 8'd117, 8'd98, 8'd79, 8'd97, 8'd158, 8'd123, 8'd122, 8'd89, 8'd127, 8'd158, 8'd122, 8'd152, 8'd98, 8'd148, 8'd156, 8'd160, 8'd87, 8'd161, 8'd87, 8'd103, 8'd148, 8'd108, 8'd85, 8'd137, 8'd151, 8'd68, 8'd72, 8'd118, 8'd99, 8'd141, 8'd125, 8'd151, 8'd147, 8'd86, 8'd104, 8'd85, 8'd84, 8'd168, 8'd114, 8'd90, 8'd79, 8'd114, 8'd112, 8'd91, 8'd157, 8'd71, 8'd70, 8'd91, 8'd128, 8'd108, 8'd133, 8'd83, 8'd89, 8'd69, 8'd51, 8'd78, 8'd112, 8'd79, 8'd81, 8'd136, 8'd110, 8'd98, 8'd95, 8'd96, 8'd175, 8'd148, 8'd140, 8'd137, 8'd123, 8'd164, 8'd96, 8'd110, 8'd96, 8'd132, 8'd125, 8'd66, 8'd123, 8'd37, 8'd121, 8'd94, 8'd107, 8'd120, 8'd129, 8'd88, 8'd149, 8'd122, 8'd108, 8'd127, 8'd76, 8'd153, 8'd94, 8'd70, 8'd108, 8'd67, 8'd84, 8'd68, 8'd144, 8'd101, 8'd97, 8'd133, 8'd154, 8'd125, 8'd66, 8'd87, 8'd117, 8'd92, 8'd76, 8'd116, 8'd112, 8'd66, 8'd91, 8'd132, 8'd96, 8'd158, 8'd98, 8'd120, 8'd94, 8'd144, 8'd145, 8'd90, 8'd159, 8'd138, 8'd83, 8'd153, 8'd105, 8'd88, 8'd120, 8'd69, 8'd65, 8'd127, 8'd82, 8'd92, 8'd91, 8'd70, 8'd92, 8'd70, 8'd143, 8'd71, 8'd119, 8'd85, 8'd154, 8'd145, 8'd115, 8'd110, 8'd118, 8'd114, 8'd92, 8'd129, 8'd135, 8'd159, 8'd129, 8'd161, 8'd90, 8'd136, 8'd75, 8'd83, 8'd158, 8'd154, 8'd119, 8'd117, 8'd93, 8'd114, 8'd92, 8'd140, 8'd115, 8'd159, 8'd104, 8'd127, 8'd159, 8'd165, 8'd149, 8'd161, 8'd110, 8'd113, 8'd166})
) cell_0_20 (
    .clk(clk),
    .input_index(index_0_19_20),
    .input_value(value_0_19_20),
    .input_result(result_0_19_20),
    .input_enable(enable_0_19_20),
    .output_index(index_0_20_21),
    .output_value(value_0_20_21),
    .output_result(result_0_20_21),
    .output_enable(enable_0_20_21)
);

wire [10-1:0] index_0_21_22;
wire [`DATA_WIDTH-1:0] value_0_21_22;
wire [`DATA_WIDTH*4:0] result_0_21_22;
wire enable_0_21_22;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd75, 8'd112, 8'd109, 8'd70, 8'd90, 8'd171, 8'd143, 8'd95, 8'd117, 8'd95, 8'd92, 8'd156, 8'd74, 8'd96, 8'd140, 8'd75, 8'd71, 8'd110, 8'd149, 8'd73, 8'd122, 8'd69, 8'd93, 8'd111, 8'd141, 8'd133, 8'd71, 8'd117, 8'd155, 8'd114, 8'd93, 8'd121, 8'd163, 8'd143, 8'd145, 8'd77, 8'd126, 8'd66, 8'd126, 8'd60, 8'd50, 8'd70, 8'd85, 8'd81, 8'd97, 8'd129, 8'd112, 8'd57, 8'd122, 8'd97, 8'd112, 8'd97, 8'd92, 8'd85, 8'd161, 8'd159, 8'd134, 8'd135, 8'd138, 8'd105, 8'd71, 8'd106, 8'd84, 8'd131, 8'd68, 8'd86, 8'd52, 8'd63, 8'd130, 8'd73, 8'd159, 8'd153, 8'd116, 8'd157, 8'd88, 8'd160, 8'd83, 8'd133, 8'd127, 8'd120, 8'd125, 8'd156, 8'd136, 8'd144, 8'd142, 8'd137, 8'd91, 8'd107, 8'd75, 8'd97, 8'd112, 8'd124, 8'd123, 8'd133, 8'd79, 8'd100, 8'd94, 8'd162, 8'd142, 8'd88, 8'd101, 8'd132, 8'd85, 8'd112, 8'd190, 8'd127, 8'd97, 8'd160, 8'd138, 8'd90, 8'd109, 8'd148, 8'd151, 8'd129, 8'd98, 8'd161, 8'd129, 8'd109, 8'd77, 8'd96, 8'd90, 8'd143, 8'd90, 8'd136, 8'd77, 8'd158, 8'd138, 8'd153, 8'd92, 8'd99, 8'd142, 8'd138, 8'd141, 8'd153, 8'd152, 8'd127, 8'd103, 8'd156, 8'd154, 8'd86, 8'd97, 8'd135, 8'd73, 8'd108, 8'd65, 8'd109, 8'd135, 8'd136, 8'd110, 8'd163, 8'd136, 8'd82, 8'd163, 8'd146, 8'd83, 8'd127, 8'd91, 8'd101, 8'd135, 8'd144, 8'd92, 8'd124, 8'd136, 8'd146, 8'd187, 8'd114, 8'd115, 8'd100, 8'd169, 8'd155, 8'd162, 8'd75, 8'd144, 8'd146, 8'd134, 8'd86, 8'd103, 8'd150, 8'd158, 8'd117, 8'd121, 8'd80, 8'd121, 8'd132, 8'd100, 8'd66, 8'd153, 8'd150, 8'd89, 8'd121, 8'd89, 8'd132, 8'd190, 8'd172, 8'd161, 8'd146, 8'd144, 8'd161, 8'd134, 8'd104, 8'd83, 8'd132, 8'd151, 8'd102, 8'd125, 8'd128, 8'd148, 8'd156, 8'd103, 8'd164, 8'd135, 8'd106, 8'd160, 8'd66, 8'd133, 8'd97, 8'd92, 8'd118, 8'd68, 8'd168, 8'd143, 8'd171, 8'd137, 8'd114, 8'd94, 8'd185, 8'd148, 8'd72, 8'd135, 8'd87, 8'd78, 8'd154, 8'd140, 8'd151, 8'd139, 8'd155, 8'd157, 8'd153, 8'd153, 8'd123, 8'd141, 8'd125, 8'd82, 8'd93, 8'd100, 8'd109, 8'd103, 8'd160, 8'd108, 8'd92, 8'd120, 8'd96, 8'd171, 8'd115, 8'd177, 8'd109, 8'd122, 8'd168, 8'd84, 8'd161, 8'd106, 8'd140, 8'd131, 8'd150, 8'd129, 8'd109, 8'd80, 8'd105, 8'd84, 8'd111, 8'd158, 8'd165, 8'd155, 8'd153, 8'd146, 8'd124, 8'd141, 8'd90, 8'd78, 8'd77, 8'd104, 8'd151, 8'd161, 8'd100, 8'd163, 8'd124, 8'd174, 8'd96, 8'd152, 8'd147, 8'd113, 8'd175, 8'd135, 8'd112, 8'd108, 8'd152, 8'd150, 8'd101, 8'd157, 8'd157, 8'd106, 8'd148, 8'd166, 8'd146, 8'd157, 8'd172, 8'd83, 8'd124, 8'd155, 8'd148, 8'd136, 8'd146, 8'd87, 8'd112, 8'd187, 8'd160, 8'd125, 8'd104, 8'd142, 8'd120, 8'd179, 8'd91, 8'd109, 8'd136, 8'd131, 8'd86, 8'd150, 8'd116, 8'd106, 8'd137, 8'd171, 8'd92, 8'd79, 8'd144, 8'd125, 8'd115, 8'd126, 8'd110, 8'd142, 8'd91, 8'd162, 8'd177, 8'd124, 8'd101, 8'd157, 8'd143, 8'd151, 8'd117, 8'd111, 8'd149, 8'd110, 8'd109, 8'd109, 8'd182, 8'd106, 8'd170, 8'd118, 8'd149, 8'd110, 8'd79, 8'd118, 8'd148, 8'd86, 8'd157, 8'd104, 8'd148, 8'd158, 8'd133, 8'd132, 8'd122, 8'd90, 8'd150, 8'd109, 8'd121, 8'd138, 8'd157, 8'd99, 8'd104, 8'd112, 8'd139, 8'd114, 8'd105, 8'd149, 8'd169, 8'd118, 8'd144, 8'd94, 8'd112, 8'd152, 8'd132, 8'd76, 8'd72, 8'd134, 8'd118, 8'd177, 8'd122, 8'd155, 8'd133, 8'd112, 8'd101, 8'd103, 8'd91, 8'd167, 8'd166, 8'd136, 8'd61, 8'd126, 8'd161, 8'd187, 8'd112, 8'd167, 8'd94, 8'd101, 8'd116, 8'd147, 8'd133, 8'd118, 8'd80, 8'd69, 8'd100, 8'd151, 8'd116, 8'd75, 8'd160, 8'd136, 8'd107, 8'd148, 8'd93, 8'd165, 8'd172, 8'd130, 8'd105, 8'd155, 8'd62, 8'd131, 8'd90, 8'd179, 8'd98, 8'd142, 8'd118, 8'd72, 8'd73, 8'd112, 8'd82, 8'd155, 8'd152, 8'd166, 8'd168, 8'd84, 8'd62, 8'd64, 8'd96, 8'd129, 8'd97, 8'd78, 8'd134, 8'd142, 8'd134, 8'd161, 8'd122, 8'd113, 8'd115, 8'd86, 8'd83, 8'd99, 8'd120, 8'd160, 8'd72, 8'd147, 8'd152, 8'd107, 8'd88, 8'd111, 8'd138, 8'd144, 8'd77, 8'd94, 8'd114, 8'd124, 8'd63, 8'd77, 8'd171, 8'd122, 8'd169, 8'd131, 8'd166, 8'd111, 8'd160, 8'd141, 8'd41, 8'd127, 8'd129, 8'd85, 8'd108, 8'd126, 8'd134, 8'd101, 8'd108, 8'd80, 8'd98, 8'd134, 8'd165, 8'd78, 8'd68, 8'd123, 8'd42, 8'd49, 8'd119, 8'd100, 8'd121, 8'd171, 8'd101, 8'd120, 8'd72, 8'd136, 8'd120, 8'd103, 8'd148, 8'd91, 8'd66, 8'd90, 8'd63, 8'd83, 8'd77, 8'd153, 8'd156, 8'd136, 8'd98, 8'd116, 8'd168, 8'd129, 8'd163, 8'd138, 8'd133, 8'd136, 8'd33, 8'd106, 8'd143, 8'd161, 8'd119, 8'd78, 8'd110, 8'd65, 8'd94, 8'd77, 8'd151, 8'd112, 8'd118, 8'd119, 8'd78, 8'd134, 8'd106, 8'd170, 8'd152, 8'd187, 8'd155, 8'd188, 8'd111, 8'd76, 8'd150, 8'd110, 8'd163, 8'd77, 8'd132, 8'd131, 8'd77, 8'd76, 8'd148, 8'd84, 8'd115, 8'd106, 8'd53, 8'd72, 8'd67, 8'd123, 8'd149, 8'd72, 8'd84, 8'd174, 8'd169, 8'd156, 8'd174, 8'd159, 8'd134, 8'd128, 8'd122, 8'd167, 8'd114, 8'd115, 8'd99, 8'd153, 8'd133, 8'd143, 8'd94, 8'd120, 8'd99, 8'd65, 8'd96, 8'd119, 8'd97, 8'd130, 8'd82, 8'd150, 8'd87, 8'd84, 8'd124, 8'd176, 8'd165, 8'd137, 8'd139, 8'd108, 8'd118, 8'd139, 8'd158, 8'd102, 8'd140, 8'd98, 8'd148, 8'd74, 8'd88, 8'd175, 8'd79, 8'd103, 8'd117, 8'd118, 8'd99, 8'd81, 8'd91, 8'd149, 8'd154, 8'd129, 8'd144, 8'd139, 8'd123, 8'd112, 8'd106, 8'd167, 8'd184, 8'd120, 8'd201, 8'd108, 8'd155, 8'd70, 8'd91, 8'd93, 8'd161, 8'd133, 8'd160, 8'd79, 8'd120, 8'd128, 8'd135, 8'd158, 8'd139, 8'd101, 8'd91, 8'd64, 8'd126, 8'd162, 8'd84, 8'd142, 8'd168, 8'd167, 8'd129, 8'd174, 8'd174, 8'd187, 8'd150, 8'd111, 8'd86, 8'd95, 8'd73, 8'd129, 8'd157, 8'd125, 8'd154, 8'd129, 8'd165, 8'd121, 8'd114, 8'd123, 8'd180, 8'd140, 8'd141, 8'd156, 8'd131, 8'd116, 8'd178, 8'd176, 8'd127, 8'd173, 8'd159, 8'd96, 8'd127, 8'd101, 8'd70, 8'd149, 8'd96, 8'd137, 8'd100, 8'd141, 8'd115, 8'd110, 8'd163, 8'd135, 8'd159, 8'd118, 8'd146, 8'd113, 8'd152, 8'd158, 8'd107, 8'd122, 8'd149, 8'd153, 8'd98, 8'd168, 8'd154, 8'd139, 8'd72, 8'd73, 8'd76, 8'd77, 8'd115, 8'd86, 8'd102, 8'd96, 8'd150, 8'd134, 8'd115, 8'd139, 8'd93, 8'd112, 8'd68, 8'd121, 8'd164, 8'd140, 8'd97, 8'd164, 8'd65, 8'd92, 8'd168, 8'd81, 8'd88, 8'd103, 8'd112, 8'd130, 8'd134, 8'd121, 8'd116, 8'd75, 8'd121, 8'd163, 8'd165, 8'd80, 8'd127, 8'd114, 8'd96, 8'd137, 8'd150, 8'd92, 8'd112, 8'd97, 8'd168, 8'd167, 8'd150, 8'd147, 8'd99, 8'd75, 8'd155, 8'd161, 8'd114, 8'd121, 8'd143, 8'd88, 8'd110, 8'd95, 8'd75, 8'd147, 8'd121, 8'd163, 8'd76, 8'd128, 8'd153})
) cell_0_21 (
    .clk(clk),
    .input_index(index_0_20_21),
    .input_value(value_0_20_21),
    .input_result(result_0_20_21),
    .input_enable(enable_0_20_21),
    .output_index(index_0_21_22),
    .output_value(value_0_21_22),
    .output_result(result_0_21_22),
    .output_enable(enable_0_21_22)
);

wire [10-1:0] index_0_22_23;
wire [`DATA_WIDTH-1:0] value_0_22_23;
wire [`DATA_WIDTH*4:0] result_0_22_23;
wire enable_0_22_23;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd114, 8'd154, 8'd116, 8'd127, 8'd104, 8'd117, 8'd127, 8'd105, 8'd150, 8'd175, 8'd199, 8'd174, 8'd126, 8'd133, 8'd112, 8'd98, 8'd91, 8'd142, 8'd96, 8'd117, 8'd99, 8'd127, 8'd176, 8'd93, 8'd71, 8'd93, 8'd115, 8'd75, 8'd117, 8'd162, 8'd117, 8'd144, 8'd124, 8'd92, 8'd138, 8'd143, 8'd166, 8'd145, 8'd174, 8'd125, 8'd114, 8'd124, 8'd149, 8'd83, 8'd117, 8'd153, 8'd137, 8'd66, 8'd81, 8'd127, 8'd136, 8'd150, 8'd135, 8'd109, 8'd150, 8'd72, 8'd114, 8'd112, 8'd158, 8'd170, 8'd85, 8'd120, 8'd86, 8'd143, 8'd120, 8'd77, 8'd116, 8'd92, 8'd123, 8'd125, 8'd112, 8'd127, 8'd105, 8'd140, 8'd157, 8'd169, 8'd117, 8'd127, 8'd161, 8'd114, 8'd100, 8'd165, 8'd162, 8'd134, 8'd140, 8'd156, 8'd80, 8'd118, 8'd85, 8'd147, 8'd93, 8'd137, 8'd94, 8'd82, 8'd119, 8'd98, 8'd164, 8'd111, 8'd122, 8'd86, 8'd175, 8'd132, 8'd150, 8'd144, 8'd83, 8'd114, 8'd168, 8'd117, 8'd188, 8'd121, 8'd144, 8'd141, 8'd106, 8'd129, 8'd139, 8'd94, 8'd59, 8'd89, 8'd103, 8'd91, 8'd133, 8'd160, 8'd120, 8'd77, 8'd164, 8'd108, 8'd124, 8'd156, 8'd94, 8'd129, 8'd126, 8'd159, 8'd138, 8'd147, 8'd121, 8'd165, 8'd154, 8'd106, 8'd157, 8'd163, 8'd77, 8'd126, 8'd143, 8'd144, 8'd140, 8'd63, 8'd65, 8'd164, 8'd153, 8'd134, 8'd85, 8'd81, 8'd86, 8'd166, 8'd166, 8'd99, 8'd117, 8'd89, 8'd102, 8'd154, 8'd98, 8'd164, 8'd130, 8'd110, 8'd123, 8'd133, 8'd165, 8'd167, 8'd121, 8'd122, 8'd82, 8'd95, 8'd135, 8'd112, 8'd164, 8'd163, 8'd113, 8'd174, 8'd135, 8'd141, 8'd161, 8'd117, 8'd159, 8'd155, 8'd116, 8'd92, 8'd171, 8'd184, 8'd115, 8'd166, 8'd76, 8'd123, 8'd198, 8'd178, 8'd165, 8'd127, 8'd148, 8'd161, 8'd136, 8'd103, 8'd133, 8'd162, 8'd145, 8'd133, 8'd104, 8'd143, 8'd121, 8'd102, 8'd113, 8'd111, 8'd186, 8'd107, 8'd144, 8'd157, 8'd179, 8'd132, 8'd87, 8'd111, 8'd88, 8'd114, 8'd146, 8'd136, 8'd150, 8'd161, 8'd82, 8'd134, 8'd163, 8'd177, 8'd177, 8'd127, 8'd178, 8'd168, 8'd133, 8'd163, 8'd98, 8'd169, 8'd168, 8'd108, 8'd111, 8'd122, 8'd117, 8'd125, 8'd182, 8'd125, 8'd166, 8'd87, 8'd160, 8'd124, 8'd125, 8'd190, 8'd137, 8'd133, 8'd117, 8'd85, 8'd123, 8'd133, 8'd141, 8'd154, 8'd127, 8'd156, 8'd114, 8'd134, 8'd160, 8'd158, 8'd69, 8'd103, 8'd177, 8'd120, 8'd122, 8'd90, 8'd70, 8'd57, 8'd124, 8'd84, 8'd155, 8'd191, 8'd188, 8'd164, 8'd104, 8'd107, 8'd166, 8'd81, 8'd163, 8'd112, 8'd187, 8'd102, 8'd173, 8'd85, 8'd178, 8'd166, 8'd100, 8'd84, 8'd138, 8'd82, 8'd115, 8'd163, 8'd74, 8'd68, 8'd110, 8'd64, 8'd53, 8'd91, 8'd135, 8'd95, 8'd120, 8'd185, 8'd163, 8'd112, 8'd119, 8'd81, 8'd119, 8'd194, 8'd141, 8'd156, 8'd168, 8'd136, 8'd96, 8'd100, 8'd85, 8'd86, 8'd75, 8'd86, 8'd169, 8'd102, 8'd88, 8'd106, 8'd103, 8'd66, 8'd76, 8'd58, 8'd89, 8'd115, 8'd165, 8'd133, 8'd96, 8'd100, 8'd68, 8'd148, 8'd92, 8'd109, 8'd106, 8'd134, 8'd93, 8'd103, 8'd157, 8'd105, 8'd89, 8'd121, 8'd113, 8'd157, 8'd142, 8'd130, 8'd77, 8'd142, 8'd83, 8'd53, 8'd69, 8'd92, 8'd63, 8'd100, 8'd100, 8'd118, 8'd83, 8'd140, 8'd70, 8'd161, 8'd95, 8'd140, 8'd158, 8'd99, 8'd58, 8'd126, 8'd84, 8'd149, 8'd113, 8'd80, 8'd77, 8'd127, 8'd135, 8'd159, 8'd73, 8'd127, 8'd122, 8'd104, 8'd66, 8'd123, 8'd74, 8'd67, 8'd77, 8'd149, 8'd172, 8'd85, 8'd116, 8'd167, 8'd132, 8'd89, 8'd74, 8'd105, 8'd131, 8'd107, 8'd128, 8'd110, 8'd54, 8'd91, 8'd80, 8'd89, 8'd147, 8'd98, 8'd91, 8'd104, 8'd93, 8'd59, 8'd87, 8'd139, 8'd145, 8'd129, 8'd147, 8'd124, 8'd118, 8'd118, 8'd118, 8'd165, 8'd113, 8'd79, 8'd98, 8'd101, 8'd96, 8'd128, 8'd85, 8'd128, 8'd61, 8'd88, 8'd94, 8'd90, 8'd93, 8'd75, 8'd117, 8'd68, 8'd85, 8'd73, 8'd119, 8'd87, 8'd77, 8'd139, 8'd137, 8'd181, 8'd149, 8'd171, 8'd130, 8'd166, 8'd171, 8'd132, 8'd109, 8'd83, 8'd77, 8'd108, 8'd61, 8'd112, 8'd92, 8'd88, 8'd122, 8'd145, 8'd176, 8'd85, 8'd98, 8'd148, 8'd132, 8'd83, 8'd102, 8'd66, 8'd121, 8'd179, 8'd152, 8'd178, 8'd101, 8'd133, 8'd125, 8'd130, 8'd150, 8'd197, 8'd181, 8'd131, 8'd69, 8'd86, 8'd89, 8'd79, 8'd134, 8'd82, 8'd183, 8'd151, 8'd175, 8'd118, 8'd89, 8'd95, 8'd92, 8'd90, 8'd151, 8'd118, 8'd124, 8'd171, 8'd113, 8'd156, 8'd98, 8'd151, 8'd157, 8'd114, 8'd214, 8'd159, 8'd94, 8'd138, 8'd84, 8'd141, 8'd156, 8'd77, 8'd98, 8'd92, 8'd157, 8'd129, 8'd114, 8'd156, 8'd134, 8'd87, 8'd149, 8'd85, 8'd134, 8'd100, 8'd112, 8'd125, 8'd146, 8'd167, 8'd105, 8'd158, 8'd168, 8'd172, 8'd170, 8'd147, 8'd182, 8'd122, 8'd92, 8'd108, 8'd141, 8'd108, 8'd83, 8'd139, 8'd142, 8'd80, 8'd158, 8'd99, 8'd128, 8'd130, 8'd72, 8'd148, 8'd112, 8'd184, 8'd110, 8'd170, 8'd100, 8'd135, 8'd183, 8'd113, 8'd131, 8'd110, 8'd189, 8'd107, 8'd167, 8'd119, 8'd163, 8'd133, 8'd136, 8'd91, 8'd144, 8'd94, 8'd69, 8'd90, 8'd165, 8'd82, 8'd90, 8'd79, 8'd138, 8'd144, 8'd109, 8'd132, 8'd162, 8'd168, 8'd183, 8'd151, 8'd99, 8'd74, 8'd117, 8'd133, 8'd123, 8'd192, 8'd139, 8'd111, 8'd137, 8'd143, 8'd82, 8'd166, 8'd81, 8'd100, 8'd136, 8'd101, 8'd133, 8'd161, 8'd83, 8'd141, 8'd116, 8'd97, 8'd147, 8'd122, 8'd140, 8'd163, 8'd116, 8'd131, 8'd122, 8'd81, 8'd171, 8'd175, 8'd185, 8'd190, 8'd94, 8'd143, 8'd146, 8'd150, 8'd127, 8'd106, 8'd134, 8'd167, 8'd97, 8'd125, 8'd112, 8'd75, 8'd109, 8'd178, 8'd97, 8'd92, 8'd123, 8'd92, 8'd128, 8'd165, 8'd129, 8'd163, 8'd161, 8'd84, 8'd135, 8'd134, 8'd97, 8'd86, 8'd156, 8'd101, 8'd188, 8'd160, 8'd114, 8'd186, 8'd115, 8'd155, 8'd178, 8'd150, 8'd114, 8'd145, 8'd156, 8'd110, 8'd115, 8'd93, 8'd170, 8'd170, 8'd112, 8'd98, 8'd170, 8'd82, 8'd80, 8'd152, 8'd145, 8'd149, 8'd155, 8'd81, 8'd164, 8'd155, 8'd190, 8'd199, 8'd173, 8'd143, 8'd174, 8'd163, 8'd206, 8'd161, 8'd192, 8'd186, 8'd143, 8'd178, 8'd186, 8'd132, 8'd128, 8'd121, 8'd134, 8'd145, 8'd166, 8'd144, 8'd94, 8'd140, 8'd145, 8'd115, 8'd115, 8'd137, 8'd100, 8'd158, 8'd149, 8'd189, 8'd169, 8'd114, 8'd183, 8'd207, 8'd120, 8'd205, 8'd167, 8'd200, 8'd190, 8'd119, 8'd157, 8'd155, 8'd191, 8'd107, 8'd104, 8'd104, 8'd151, 8'd107, 8'd109, 8'd153, 8'd120, 8'd96, 8'd112, 8'd84, 8'd85, 8'd121, 8'd169, 8'd107, 8'd103, 8'd119, 8'd112, 8'd162, 8'd182, 8'd177, 8'd132, 8'd145, 8'd110, 8'd176, 8'd178, 8'd142, 8'd184, 8'd123, 8'd164, 8'd109, 8'd114, 8'd110, 8'd81, 8'd157, 8'd114, 8'd112, 8'd149, 8'd105, 8'd142, 8'd162, 8'd90, 8'd168, 8'd79, 8'd131, 8'd116, 8'd145, 8'd76, 8'd148, 8'd139, 8'd166, 8'd101, 8'd99, 8'd111, 8'd167, 8'd72, 8'd139, 8'd161, 8'd169, 8'd155, 8'd98, 8'd143, 8'd158})
) cell_0_22 (
    .clk(clk),
    .input_index(index_0_21_22),
    .input_value(value_0_21_22),
    .input_result(result_0_21_22),
    .input_enable(enable_0_21_22),
    .output_index(index_0_22_23),
    .output_value(value_0_22_23),
    .output_result(result_0_22_23),
    .output_enable(enable_0_22_23)
);

wire [10-1:0] index_0_23_24;
wire [`DATA_WIDTH-1:0] value_0_23_24;
wire [`DATA_WIDTH*4:0] result_0_23_24;
wire enable_0_23_24;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd76, 8'd115, 8'd164, 8'd167, 8'd148, 8'd124, 8'd116, 8'd118, 8'd53, 8'd65, 8'd47, 8'd84, 8'd116, 8'd113, 8'd50, 8'd94, 8'd151, 8'd80, 8'd117, 8'd122, 8'd79, 8'd160, 8'd117, 8'd144, 8'd140, 8'd73, 8'd129, 8'd97, 8'd82, 8'd154, 8'd101, 8'd146, 8'd117, 8'd114, 8'd116, 8'd158, 8'd149, 8'd118, 8'd144, 8'd142, 8'd126, 8'd122, 8'd78, 8'd128, 8'd130, 8'd88, 8'd82, 8'd129, 8'd160, 8'd97, 8'd121, 8'd133, 8'd147, 8'd137, 8'd110, 8'd110, 8'd99, 8'd98, 8'd102, 8'd96, 8'd150, 8'd93, 8'd97, 8'd169, 8'd163, 8'd167, 8'd157, 8'd125, 8'd184, 8'd103, 8'd108, 8'd148, 8'd155, 8'd166, 8'd167, 8'd160, 8'd139, 8'd77, 8'd119, 8'd66, 8'd92, 8'd113, 8'd128, 8'd98, 8'd93, 8'd78, 8'd124, 8'd160, 8'd198, 8'd185, 8'd120, 8'd171, 8'd130, 8'd119, 8'd83, 8'd135, 8'd109, 8'd124, 8'd104, 8'd119, 8'd119, 8'd163, 8'd153, 8'd94, 8'd90, 8'd145, 8'd126, 8'd113, 8'd149, 8'd137, 8'd158, 8'd97, 8'd141, 8'd100, 8'd101, 8'd198, 8'd130, 8'd168, 8'd163, 8'd160, 8'd101, 8'd158, 8'd93, 8'd105, 8'd128, 8'd118, 8'd126, 8'd172, 8'd109, 8'd112, 8'd121, 8'd121, 8'd82, 8'd85, 8'd128, 8'd87, 8'd174, 8'd149, 8'd84, 8'd123, 8'd109, 8'd100, 8'd157, 8'd149, 8'd145, 8'd180, 8'd110, 8'd149, 8'd91, 8'd155, 8'd136, 8'd101, 8'd158, 8'd78, 8'd82, 8'd102, 8'd95, 8'd97, 8'd162, 8'd161, 8'd178, 8'd86, 8'd117, 8'd155, 8'd130, 8'd80, 8'd123, 8'd95, 8'd144, 8'd161, 8'd181, 8'd160, 8'd126, 8'd188, 8'd124, 8'd112, 8'd93, 8'd134, 8'd86, 8'd67, 8'd72, 8'd121, 8'd69, 8'd135, 8'd158, 8'd72, 8'd97, 8'd180, 8'd172, 8'd186, 8'd121, 8'd163, 8'd175, 8'd159, 8'd120, 8'd92, 8'd152, 8'd75, 8'd179, 8'd194, 8'd176, 8'd130, 8'd117, 8'd162, 8'd131, 8'd105, 8'd84, 8'd147, 8'd150, 8'd140, 8'd89, 8'd150, 8'd69, 8'd120, 8'd145, 8'd167, 8'd130, 8'd159, 8'd105, 8'd99, 8'd168, 8'd92, 8'd119, 8'd159, 8'd122, 8'd127, 8'd186, 8'd103, 8'd167, 8'd109, 8'd112, 8'd180, 8'd164, 8'd144, 8'd136, 8'd162, 8'd67, 8'd92, 8'd102, 8'd119, 8'd121, 8'd135, 8'd175, 8'd190, 8'd186, 8'd141, 8'd114, 8'd108, 8'd118, 8'd147, 8'd138, 8'd132, 8'd172, 8'd174, 8'd173, 8'd126, 8'd99, 8'd135, 8'd85, 8'd143, 8'd137, 8'd94, 8'd90, 8'd125, 8'd82, 8'd154, 8'd88, 8'd121, 8'd108, 8'd79, 8'd133, 8'd136, 8'd108, 8'd136, 8'd131, 8'd109, 8'd144, 8'd83, 8'd144, 8'd129, 8'd133, 8'd152, 8'd181, 8'd96, 8'd119, 8'd108, 8'd70, 8'd141, 8'd97, 8'd78, 8'd162, 8'd131, 8'd102, 8'd86, 8'd71, 8'd71, 8'd160, 8'd116, 8'd79, 8'd120, 8'd100, 8'd131, 8'd90, 8'd173, 8'd103, 8'd139, 8'd102, 8'd90, 8'd133, 8'd201, 8'd171, 8'd105, 8'd114, 8'd115, 8'd97, 8'd101, 8'd152, 8'd98, 8'd166, 8'd159, 8'd121, 8'd57, 8'd109, 8'd167, 8'd163, 8'd149, 8'd112, 8'd133, 8'd102, 8'd80, 8'd112, 8'd143, 8'd143, 8'd92, 8'd159, 8'd152, 8'd184, 8'd123, 8'd102, 8'd93, 8'd96, 8'd126, 8'd76, 8'd95, 8'd134, 8'd148, 8'd80, 8'd128, 8'd63, 8'd141, 8'd109, 8'd96, 8'd152, 8'd141, 8'd70, 8'd70, 8'd65, 8'd83, 8'd155, 8'd125, 8'd80, 8'd109, 8'd151, 8'd93, 8'd101, 8'd127, 8'd155, 8'd89, 8'd63, 8'd103, 8'd76, 8'd143, 8'd152, 8'd122, 8'd107, 8'd65, 8'd101, 8'd83, 8'd91, 8'd182, 8'd136, 8'd149, 8'd151, 8'd83, 8'd112, 8'd132, 8'd85, 8'd148, 8'd127, 8'd54, 8'd71, 8'd144, 8'd126, 8'd110, 8'd130, 8'd97, 8'd38, 8'd104, 8'd87, 8'd79, 8'd89, 8'd79, 8'd167, 8'd132, 8'd86, 8'd114, 8'd157, 8'd107, 8'd163, 8'd125, 8'd113, 8'd72, 8'd113, 8'd62, 8'd136, 8'd70, 8'd148, 8'd53, 8'd127, 8'd90, 8'd85, 8'd106, 8'd137, 8'd83, 8'd61, 8'd111, 8'd79, 8'd114, 8'd127, 8'd142, 8'd118, 8'd83, 8'd146, 8'd76, 8'd96, 8'd121, 8'd109, 8'd89, 8'd142, 8'd66, 8'd122, 8'd108, 8'd172, 8'd103, 8'd83, 8'd109, 8'd72, 8'd137, 8'd78, 8'd197, 8'd217, 8'd109, 8'd125, 8'd96, 8'd100, 8'd130, 8'd130, 8'd156, 8'd134, 8'd134, 8'd86, 8'd136, 8'd82, 8'd144, 8'd137, 8'd153, 8'd134, 8'd96, 8'd163, 8'd138, 8'd140, 8'd109, 8'd69, 8'd138, 8'd61, 8'd144, 8'd118, 8'd190, 8'd184, 8'd119, 8'd115, 8'd92, 8'd94, 8'd115, 8'd100, 8'd156, 8'd118, 8'd101, 8'd150, 8'd98, 8'd153, 8'd125, 8'd169, 8'd127, 8'd165, 8'd110, 8'd154, 8'd130, 8'd161, 8'd95, 8'd151, 8'd107, 8'd65, 8'd133, 8'd90, 8'd145, 8'd223, 8'd131, 8'd137, 8'd143, 8'd82, 8'd125, 8'd129, 8'd112, 8'd113, 8'd77, 8'd131, 8'd106, 8'd101, 8'd83, 8'd164, 8'd133, 8'd144, 8'd97, 8'd167, 8'd151, 8'd137, 8'd109, 8'd142, 8'd95, 8'd72, 8'd80, 8'd141, 8'd119, 8'd122, 8'd148, 8'd109, 8'd165, 8'd106, 8'd170, 8'd104, 8'd147, 8'd96, 8'd115, 8'd162, 8'd125, 8'd86, 8'd77, 8'd98, 8'd102, 8'd85, 8'd122, 8'd115, 8'd111, 8'd66, 8'd83, 8'd88, 8'd121, 8'd135, 8'd138, 8'd91, 8'd155, 8'd172, 8'd97, 8'd147, 8'd157, 8'd144, 8'd105, 8'd106, 8'd118, 8'd134, 8'd166, 8'd154, 8'd121, 8'd91, 8'd151, 8'd134, 8'd143, 8'd180, 8'd165, 8'd91, 8'd121, 8'd144, 8'd51, 8'd82, 8'd119, 8'd99, 8'd122, 8'd165, 8'd97, 8'd127, 8'd95, 8'd103, 8'd103, 8'd77, 8'd71, 8'd130, 8'd179, 8'd138, 8'd150, 8'd154, 8'd154, 8'd181, 8'd153, 8'd175, 8'd121, 8'd134, 8'd159, 8'd145, 8'd78, 8'd116, 8'd93, 8'd105, 8'd125, 8'd138, 8'd103, 8'd155, 8'd105, 8'd126, 8'd116, 8'd101, 8'd62, 8'd132, 8'd135, 8'd114, 8'd81, 8'd111, 8'd100, 8'd143, 8'd115, 8'd180, 8'd144, 8'd130, 8'd127, 8'd163, 8'd115, 8'd84, 8'd121, 8'd82, 8'd89, 8'd130, 8'd80, 8'd111, 8'd75, 8'd99, 8'd113, 8'd89, 8'd145, 8'd139, 8'd63, 8'd95, 8'd118, 8'd77, 8'd127, 8'd101, 8'd156, 8'd147, 8'd79, 8'd91, 8'd160, 8'd151, 8'd167, 8'd137, 8'd125, 8'd81, 8'd128, 8'd67, 8'd138, 8'd91, 8'd94, 8'd142, 8'd133, 8'd137, 8'd102, 8'd83, 8'd131, 8'd104, 8'd62, 8'd62, 8'd122, 8'd131, 8'd64, 8'd72, 8'd110, 8'd97, 8'd136, 8'd94, 8'd91, 8'd148, 8'd114, 8'd137, 8'd75, 8'd152, 8'd141, 8'd132, 8'd116, 8'd82, 8'd125, 8'd154, 8'd96, 8'd83, 8'd132, 8'd118, 8'd154, 8'd90, 8'd81, 8'd123, 8'd102, 8'd133, 8'd106, 8'd91, 8'd102, 8'd126, 8'd43, 8'd131, 8'd59, 8'd141, 8'd96, 8'd77, 8'd53, 8'd102, 8'd88, 8'd132, 8'd115, 8'd127, 8'd152, 8'd145, 8'd120, 8'd108, 8'd74, 8'd163, 8'd153, 8'd156, 8'd128, 8'd154, 8'd147, 8'd79, 8'd54, 8'd105, 8'd132, 8'd141, 8'd105, 8'd53, 8'd73, 8'd103, 8'd77, 8'd62, 8'd133, 8'd73, 8'd92, 8'd132, 8'd166, 8'd137, 8'd96, 8'd80, 8'd126, 8'd134, 8'd74, 8'd99, 8'd147, 8'd153, 8'd161, 8'd84, 8'd81, 8'd99, 8'd162, 8'd105, 8'd119, 8'd114, 8'd146, 8'd123, 8'd99, 8'd70, 8'd124, 8'd111, 8'd111, 8'd93, 8'd157, 8'd72, 8'd86, 8'd146, 8'd76, 8'd130, 8'd114})
) cell_0_23 (
    .clk(clk),
    .input_index(index_0_22_23),
    .input_value(value_0_22_23),
    .input_result(result_0_22_23),
    .input_enable(enable_0_22_23),
    .output_index(index_0_23_24),
    .output_value(value_0_23_24),
    .output_result(result_0_23_24),
    .output_enable(enable_0_23_24)
);

wire [10-1:0] index_0_24_25;
wire [`DATA_WIDTH-1:0] value_0_24_25;
wire [`DATA_WIDTH*4:0] result_0_24_25;
wire enable_0_24_25;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd157, 8'd120, 8'd131, 8'd83, 8'd103, 8'd135, 8'd117, 8'd105, 8'd152, 8'd151, 8'd187, 8'd181, 8'd174, 8'd187, 8'd144, 8'd83, 8'd116, 8'd113, 8'd94, 8'd106, 8'd139, 8'd127, 8'd150, 8'd123, 8'd145, 8'd127, 8'd113, 8'd116, 8'd85, 8'd134, 8'd78, 8'd127, 8'd140, 8'd73, 8'd120, 8'd91, 8'd113, 8'd161, 8'd156, 8'd111, 8'd92, 8'd123, 8'd159, 8'd143, 8'd71, 8'd105, 8'd169, 8'd169, 8'd186, 8'd169, 8'd136, 8'd175, 8'd150, 8'd74, 8'd70, 8'd91, 8'd112, 8'd167, 8'd142, 8'd127, 8'd97, 8'd63, 8'd158, 8'd76, 8'd142, 8'd63, 8'd93, 8'd117, 8'd78, 8'd120, 8'd126, 8'd121, 8'd148, 8'd121, 8'd72, 8'd176, 8'd94, 8'd134, 8'd112, 8'd138, 8'd136, 8'd82, 8'd158, 8'd104, 8'd81, 8'd150, 8'd133, 8'd148, 8'd85, 8'd158, 8'd120, 8'd94, 8'd107, 8'd107, 8'd98, 8'd61, 8'd103, 8'd70, 8'd42, 8'd105, 8'd126, 8'd112, 8'd119, 8'd150, 8'd177, 8'd140, 8'd188, 8'd167, 8'd76, 8'd80, 8'd132, 8'd141, 8'd71, 8'd87, 8'd135, 8'd156, 8'd75, 8'd75, 8'd126, 8'd87, 8'd131, 8'd150, 8'd158, 8'd90, 8'd114, 8'd52, 8'd57, 8'd100, 8'd114, 8'd37, 8'd49, 8'd67, 8'd142, 8'd112, 8'd109, 8'd164, 8'd83, 8'd91, 8'd165, 8'd122, 8'd71, 8'd100, 8'd98, 8'd76, 8'd74, 8'd103, 8'd81, 8'd133, 8'd95, 8'd83, 8'd147, 8'd126, 8'd80, 8'd74, 8'd111, 8'd103, 8'd133, 8'd104, 8'd130, 8'd148, 8'd65, 8'd131, 8'd84, 8'd97, 8'd158, 8'd175, 8'd103, 8'd160, 8'd141, 8'd107, 8'd77, 8'd98, 8'd83, 8'd93, 8'd118, 8'd92, 8'd84, 8'd175, 8'd105, 8'd89, 8'd101, 8'd181, 8'd174, 8'd94, 8'd153, 8'd89, 8'd64, 8'd118, 8'd115, 8'd117, 8'd50, 8'd129, 8'd89, 8'd113, 8'd121, 8'd79, 8'd77, 8'd88, 8'd157, 8'd93, 8'd105, 8'd133, 8'd125, 8'd80, 8'd100, 8'd154, 8'd166, 8'd134, 8'd115, 8'd117, 8'd147, 8'd172, 8'd112, 8'd168, 8'd150, 8'd145, 8'd120, 8'd76, 8'd71, 8'd77, 8'd166, 8'd69, 8'd138, 8'd104, 8'd95, 8'd152, 8'd117, 8'd154, 8'd73, 8'd152, 8'd162, 8'd162, 8'd119, 8'd159, 8'd97, 8'd94, 8'd163, 8'd104, 8'd182, 8'd143, 8'd175, 8'd138, 8'd85, 8'd74, 8'd65, 8'd96, 8'd51, 8'd115, 8'd91, 8'd107, 8'd146, 8'd102, 8'd96, 8'd121, 8'd117, 8'd101, 8'd148, 8'd137, 8'd87, 8'd150, 8'd85, 8'd153, 8'd82, 8'd150, 8'd128, 8'd106, 8'd185, 8'd194, 8'd172, 8'd132, 8'd164, 8'd120, 8'd145, 8'd130, 8'd102, 8'd138, 8'd170, 8'd171, 8'd103, 8'd120, 8'd88, 8'd103, 8'd155, 8'd130, 8'd156, 8'd132, 8'd87, 8'd104, 8'd153, 8'd127, 8'd152, 8'd110, 8'd167, 8'd190, 8'd144, 8'd116, 8'd144, 8'd128, 8'd128, 8'd123, 8'd72, 8'd72, 8'd51, 8'd113, 8'd98, 8'd111, 8'd123, 8'd71, 8'd97, 8'd140, 8'd116, 8'd113, 8'd87, 8'd93, 8'd168, 8'd99, 8'd111, 8'd121, 8'd154, 8'd101, 8'd195, 8'd116, 8'd160, 8'd126, 8'd170, 8'd156, 8'd108, 8'd154, 8'd93, 8'd138, 8'd105, 8'd71, 8'd78, 8'd138, 8'd87, 8'd163, 8'd165, 8'd116, 8'd162, 8'd142, 8'd129, 8'd80, 8'd127, 8'd166, 8'd117, 8'd160, 8'd142, 8'd160, 8'd191, 8'd177, 8'd187, 8'd100, 8'd130, 8'd112, 8'd130, 8'd139, 8'd169, 8'd100, 8'd148, 8'd82, 8'd155, 8'd127, 8'd130, 8'd101, 8'd140, 8'd113, 8'd101, 8'd130, 8'd111, 8'd118, 8'd117, 8'd80, 8'd129, 8'd106, 8'd160, 8'd127, 8'd213, 8'd121, 8'd153, 8'd72, 8'd106, 8'd101, 8'd80, 8'd142, 8'd162, 8'd104, 8'd131, 8'd129, 8'd164, 8'd137, 8'd153, 8'd95, 8'd136, 8'd83, 8'd139, 8'd170, 8'd100, 8'd142, 8'd112, 8'd132, 8'd90, 8'd75, 8'd102, 8'd174, 8'd124, 8'd168, 8'd151, 8'd83, 8'd79, 8'd146, 8'd92, 8'd96, 8'd158, 8'd85, 8'd83, 8'd79, 8'd162, 8'd168, 8'd166, 8'd130, 8'd137, 8'd98, 8'd81, 8'd117, 8'd169, 8'd160, 8'd127, 8'd69, 8'd90, 8'd109, 8'd72, 8'd108, 8'd116, 8'd144, 8'd71, 8'd96, 8'd154, 8'd70, 8'd152, 8'd103, 8'd88, 8'd144, 8'd113, 8'd109, 8'd97, 8'd91, 8'd139, 8'd148, 8'd128, 8'd43, 8'd85, 8'd44, 8'd148, 8'd159, 8'd66, 8'd89, 8'd74, 8'd81, 8'd96, 8'd118, 8'd114, 8'd168, 8'd151, 8'd84, 8'd148, 8'd114, 8'd60, 8'd68, 8'd148, 8'd113, 8'd93, 8'd93, 8'd172, 8'd168, 8'd86, 8'd119, 8'd120, 8'd88, 8'd39, 8'd78, 8'd86, 8'd105, 8'd136, 8'd93, 8'd113, 8'd84, 8'd148, 8'd164, 8'd107, 8'd124, 8'd95, 8'd127, 8'd85, 8'd55, 8'd140, 8'd137, 8'd105, 8'd62, 8'd122, 8'd116, 8'd113, 8'd114, 8'd130, 8'd146, 8'd76, 8'd108, 8'd76, 8'd61, 8'd18, 8'd39, 8'd68, 8'd95, 8'd45, 8'd44, 8'd128, 8'd83, 8'd89, 8'd172, 8'd64, 8'd118, 8'd56, 8'd108, 8'd63, 8'd121, 8'd80, 8'd139, 8'd147, 8'd147, 8'd88, 8'd147, 8'd132, 8'd74, 8'd146, 8'd126, 8'd69, 8'd88, 8'd67, 8'd132, 8'd85, 8'd84, 8'd118, 8'd48, 8'd123, 8'd63, 8'd164, 8'd156, 8'd104, 8'd88, 8'd119, 8'd71, 8'd134, 8'd140, 8'd74, 8'd95, 8'd74, 8'd142, 8'd123, 8'd145, 8'd132, 8'd130, 8'd149, 8'd82, 8'd101, 8'd50, 8'd56, 8'd78, 8'd59, 8'd122, 8'd111, 8'd115, 8'd55, 8'd101, 8'd86, 8'd75, 8'd140, 8'd65, 8'd61, 8'd75, 8'd118, 8'd137, 8'd121, 8'd83, 8'd101, 8'd148, 8'd88, 8'd161, 8'd172, 8'd75, 8'd99, 8'd122, 8'd57, 8'd125, 8'd110, 8'd60, 8'd69, 8'd81, 8'd94, 8'd112, 8'd67, 8'd140, 8'd143, 8'd62, 8'd87, 8'd125, 8'd111, 8'd75, 8'd75, 8'd98, 8'd115, 8'd115, 8'd106, 8'd179, 8'd165, 8'd103, 8'd104, 8'd110, 8'd120, 8'd68, 8'd75, 8'd139, 8'd93, 8'd151, 8'd169, 8'd89, 8'd117, 8'd147, 8'd84, 8'd60, 8'd159, 8'd105, 8'd139, 8'd101, 8'd125, 8'd160, 8'd145, 8'd153, 8'd102, 8'd120, 8'd141, 8'd175, 8'd114, 8'd103, 8'd113, 8'd110, 8'd133, 8'd76, 8'd129, 8'd85, 8'd111, 8'd145, 8'd118, 8'd134, 8'd123, 8'd163, 8'd97, 8'd164, 8'd129, 8'd161, 8'd96, 8'd151, 8'd155, 8'd111, 8'd129, 8'd103, 8'd177, 8'd100, 8'd156, 8'd160, 8'd70, 8'd153, 8'd165, 8'd146, 8'd132, 8'd108, 8'd154, 8'd188, 8'd138, 8'd135, 8'd150, 8'd138, 8'd170, 8'd146, 8'd155, 8'd122, 8'd144, 8'd126, 8'd182, 8'd151, 8'd125, 8'd192, 8'd111, 8'd125, 8'd113, 8'd110, 8'd155, 8'd126, 8'd89, 8'd126, 8'd130, 8'd144, 8'd167, 8'd137, 8'd129, 8'd99, 8'd109, 8'd109, 8'd126, 8'd112, 8'd165, 8'd123, 8'd126, 8'd150, 8'd216, 8'd188, 8'd126, 8'd159, 8'd143, 8'd155, 8'd162, 8'd164, 8'd110, 8'd146, 8'd178, 8'd74, 8'd94, 8'd137, 8'd148, 8'd97, 8'd125, 8'd114, 8'd99, 8'd157, 8'd113, 8'd179, 8'd126, 8'd135, 8'd167, 8'd128, 8'd132, 8'd155, 8'd138, 8'd138, 8'd174, 8'd153, 8'd172, 8'd186, 8'd98, 8'd159, 8'd107, 8'd123, 8'd162, 8'd82, 8'd100, 8'd113, 8'd90, 8'd140, 8'd142, 8'd106, 8'd120, 8'd167, 8'd88, 8'd109, 8'd141, 8'd120, 8'd158, 8'd78, 8'd142, 8'd126, 8'd163, 8'd69, 8'd103, 8'd158, 8'd120, 8'd71, 8'd76, 8'd97, 8'd156, 8'd128, 8'd117, 8'd111, 8'd70, 8'd165, 8'd81, 8'd148})
) cell_0_24 (
    .clk(clk),
    .input_index(index_0_23_24),
    .input_value(value_0_23_24),
    .input_result(result_0_23_24),
    .input_enable(enable_0_23_24),
    .output_index(index_0_24_25),
    .output_value(value_0_24_25),
    .output_result(result_0_24_25),
    .output_enable(enable_0_24_25)
);

wire [10-1:0] index_0_25_26;
wire [`DATA_WIDTH-1:0] value_0_25_26;
wire [`DATA_WIDTH*4:0] result_0_25_26;
wire enable_0_25_26;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd120, 8'd91, 8'd169, 8'd108, 8'd120, 8'd156, 8'd64, 8'd158, 8'd116, 8'd121, 8'd48, 8'd69, 8'd117, 8'd60, 8'd49, 8'd91, 8'd96, 8'd153, 8'd93, 8'd114, 8'd169, 8'd92, 8'd159, 8'd80, 8'd146, 8'd108, 8'd109, 8'd91, 8'd109, 8'd124, 8'd111, 8'd120, 8'd73, 8'd147, 8'd169, 8'd99, 8'd66, 8'd157, 8'd132, 8'd102, 8'd102, 8'd68, 8'd65, 8'd72, 8'd137, 8'd107, 8'd120, 8'd78, 8'd130, 8'd154, 8'd148, 8'd121, 8'd132, 8'd83, 8'd160, 8'd129, 8'd120, 8'd159, 8'd107, 8'd152, 8'd171, 8'd137, 8'd143, 8'd184, 8'd113, 8'd78, 8'd153, 8'd144, 8'd85, 8'd109, 8'd81, 8'd130, 8'd43, 8'd75, 8'd66, 8'd48, 8'd33, 8'd107, 8'd127, 8'd64, 8'd73, 8'd157, 8'd77, 8'd74, 8'd111, 8'd89, 8'd133, 8'd114, 8'd157, 8'd164, 8'd123, 8'd88, 8'd97, 8'd136, 8'd138, 8'd171, 8'd85, 8'd108, 8'd113, 8'd88, 8'd106, 8'd125, 8'd105, 8'd90, 8'd57, 8'd48, 8'd101, 8'd46, 8'd103, 8'd170, 8'd150, 8'd144, 8'd120, 8'd174, 8'd72, 8'd88, 8'd164, 8'd136, 8'd69, 8'd111, 8'd128, 8'd156, 8'd176, 8'd180, 8'd127, 8'd166, 8'd113, 8'd175, 8'd101, 8'd129, 8'd116, 8'd158, 8'd104, 8'd150, 8'd123, 8'd82, 8'd108, 8'd127, 8'd86, 8'd132, 8'd104, 8'd177, 8'd141, 8'd56, 8'd131, 8'd156, 8'd127, 8'd112, 8'd86, 8'd92, 8'd128, 8'd99, 8'd120, 8'd94, 8'd102, 8'd125, 8'd147, 8'd164, 8'd116, 8'd99, 8'd166, 8'd80, 8'd141, 8'd78, 8'd88, 8'd151, 8'd139, 8'd99, 8'd90, 8'd112, 8'd89, 8'd56, 8'd137, 8'd128, 8'd105, 8'd99, 8'd119, 8'd128, 8'd106, 8'd80, 8'd108, 8'd110, 8'd111, 8'd148, 8'd88, 8'd170, 8'd95, 8'd77, 8'd179, 8'd102, 8'd143, 8'd145, 8'd59, 8'd131, 8'd95, 8'd106, 8'd166, 8'd61, 8'd52, 8'd121, 8'd104, 8'd140, 8'd83, 8'd97, 8'd126, 8'd127, 8'd120, 8'd121, 8'd130, 8'd110, 8'd129, 8'd110, 8'd100, 8'd156, 8'd114, 8'd179, 8'd128, 8'd103, 8'd121, 8'd122, 8'd135, 8'd152, 8'd70, 8'd112, 8'd67, 8'd129, 8'd68, 8'd123, 8'd98, 8'd155, 8'd80, 8'd167, 8'd86, 8'd166, 8'd116, 8'd138, 8'd122, 8'd67, 8'd156, 8'd104, 8'd157, 8'd136, 8'd176, 8'd104, 8'd114, 8'd85, 8'd114, 8'd57, 8'd87, 8'd164, 8'd115, 8'd102, 8'd150, 8'd53, 8'd86, 8'd84, 8'd127, 8'd162, 8'd118, 8'd103, 8'd103, 8'd78, 8'd142, 8'd84, 8'd141, 8'd94, 8'd150, 8'd153, 8'd111, 8'd140, 8'd116, 8'd140, 8'd119, 8'd160, 8'd84, 8'd87, 8'd144, 8'd170, 8'd118, 8'd88, 8'd132, 8'd116, 8'd50, 8'd64, 8'd103, 8'd82, 8'd148, 8'd124, 8'd92, 8'd54, 8'd70, 8'd57, 8'd89, 8'd130, 8'd173, 8'd108, 8'd166, 8'd86, 8'd121, 8'd81, 8'd68, 8'd92, 8'd118, 8'd140, 8'd91, 8'd104, 8'd147, 8'd115, 8'd103, 8'd53, 8'd65, 8'd151, 8'd105, 8'd147, 8'd62, 8'd59, 8'd87, 8'd40, 8'd68, 8'd124, 8'd88, 8'd132, 8'd128, 8'd161, 8'd148, 8'd155, 8'd71, 8'd85, 8'd126, 8'd84, 8'd101, 8'd114, 8'd153, 8'd92, 8'd147, 8'd121, 8'd128, 8'd63, 8'd61, 8'd86, 8'd64, 8'd133, 8'd115, 8'd93, 8'd52, 8'd129, 8'd115, 8'd111, 8'd128, 8'd145, 8'd128, 8'd109, 8'd80, 8'd161, 8'd151, 8'd123, 8'd107, 8'd65, 8'd90, 8'd100, 8'd92, 8'd76, 8'd167, 8'd165, 8'd146, 8'd83, 8'd121, 8'd107, 8'd117, 8'd126, 8'd69, 8'd124, 8'd51, 8'd106, 8'd91, 8'd68, 8'd169, 8'd151, 8'd157, 8'd121, 8'd127, 8'd134, 8'd149, 8'd117, 8'd89, 8'd65, 8'd63, 8'd125, 8'd146, 8'd58, 8'd110, 8'd88, 8'd91, 8'd102, 8'd62, 8'd156, 8'd170, 8'd111, 8'd90, 8'd105, 8'd134, 8'd80, 8'd116, 8'd167, 8'd124, 8'd139, 8'd203, 8'd159, 8'd135, 8'd130, 8'd164, 8'd118, 8'd171, 8'd179, 8'd146, 8'd144, 8'd79, 8'd76, 8'd79, 8'd91, 8'd83, 8'd113, 8'd113, 8'd173, 8'd130, 8'd166, 8'd114, 8'd148, 8'd88, 8'd122, 8'd103, 8'd95, 8'd94, 8'd207, 8'd155, 8'd123, 8'd117, 8'd178, 8'd149, 8'd97, 8'd143, 8'd171, 8'd176, 8'd94, 8'd126, 8'd80, 8'd122, 8'd142, 8'd91, 8'd190, 8'd174, 8'd152, 8'd178, 8'd119, 8'd112, 8'd142, 8'd85, 8'd134, 8'd73, 8'd85, 8'd109, 8'd200, 8'd179, 8'd196, 8'd124, 8'd112, 8'd180, 8'd115, 8'd108, 8'd189, 8'd139, 8'd130, 8'd62, 8'd115, 8'd112, 8'd145, 8'd142, 8'd115, 8'd204, 8'd214, 8'd188, 8'd151, 8'd145, 8'd94, 8'd128, 8'd137, 8'd106, 8'd75, 8'd91, 8'd102, 8'd176, 8'd181, 8'd112, 8'd101, 8'd171, 8'd145, 8'd179, 8'd158, 8'd105, 8'd123, 8'd58, 8'd42, 8'd97, 8'd146, 8'd158, 8'd118, 8'd208, 8'd216, 8'd138, 8'd139, 8'd137, 8'd68, 8'd98, 8'd106, 8'd121, 8'd116, 8'd44, 8'd65, 8'd147, 8'd75, 8'd76, 8'd166, 8'd123, 8'd76, 8'd101, 8'd123, 8'd146, 8'd100, 8'd102, 8'd72, 8'd112, 8'd154, 8'd141, 8'd131, 8'd134, 8'd221, 8'd113, 8'd175, 8'd164, 8'd85, 8'd81, 8'd166, 8'd63, 8'd57, 8'd48, 8'd92, 8'd140, 8'd117, 8'd75, 8'd104, 8'd152, 8'd78, 8'd147, 8'd72, 8'd139, 8'd47, 8'd130, 8'd88, 8'd92, 8'd116, 8'd93, 8'd136, 8'd185, 8'd151, 8'd172, 8'd95, 8'd139, 8'd93, 8'd138, 8'd97, 8'd127, 8'd145, 8'd100, 8'd50, 8'd89, 8'd147, 8'd80, 8'd99, 8'd123, 8'd139, 8'd131, 8'd59, 8'd117, 8'd64, 8'd104, 8'd107, 8'd101, 8'd125, 8'd91, 8'd157, 8'd138, 8'd206, 8'd193, 8'd180, 8'd121, 8'd161, 8'd97, 8'd169, 8'd118, 8'd104, 8'd158, 8'd116, 8'd130, 8'd151, 8'd145, 8'd124, 8'd127, 8'd78, 8'd141, 8'd144, 8'd92, 8'd122, 8'd131, 8'd148, 8'd157, 8'd150, 8'd108, 8'd179, 8'd126, 8'd143, 8'd135, 8'd151, 8'd110, 8'd116, 8'd121, 8'd133, 8'd104, 8'd140, 8'd126, 8'd96, 8'd139, 8'd143, 8'd86, 8'd97, 8'd61, 8'd111, 8'd93, 8'd81, 8'd100, 8'd91, 8'd159, 8'd163, 8'd134, 8'd162, 8'd130, 8'd156, 8'd112, 8'd142, 8'd176, 8'd119, 8'd154, 8'd97, 8'd133, 8'd86, 8'd102, 8'd138, 8'd164, 8'd152, 8'd126, 8'd119, 8'd157, 8'd83, 8'd110, 8'd114, 8'd129, 8'd94, 8'd73, 8'd147, 8'd169, 8'd94, 8'd131, 8'd143, 8'd158, 8'd69, 8'd150, 8'd155, 8'd145, 8'd121, 8'd78, 8'd139, 8'd155, 8'd141, 8'd82, 8'd120, 8'd113, 8'd73, 8'd140, 8'd106, 8'd109, 8'd69, 8'd129, 8'd165, 8'd152, 8'd148, 8'd104, 8'd97, 8'd179, 8'd81, 8'd167, 8'd136, 8'd128, 8'd99, 8'd98, 8'd134, 8'd152, 8'd119, 8'd102, 8'd90, 8'd169, 8'd88, 8'd139, 8'd117, 8'd132, 8'd84, 8'd124, 8'd178, 8'd138, 8'd140, 8'd155, 8'd170, 8'd186, 8'd112, 8'd108, 8'd92, 8'd95, 8'd102, 8'd89, 8'd99, 8'd144, 8'd109, 8'd81, 8'd83, 8'd132, 8'd155, 8'd116, 8'd122, 8'd112, 8'd109, 8'd157, 8'd165, 8'd148, 8'd119, 8'd129, 8'd123, 8'd117, 8'd183, 8'd160, 8'd138, 8'd131, 8'd140, 8'd136, 8'd84, 8'd153, 8'd153, 8'd143, 8'd128, 8'd115, 8'd92, 8'd157, 8'd160, 8'd135, 8'd112, 8'd151, 8'd77, 8'd113, 8'd100, 8'd78, 8'd157, 8'd154, 8'd101, 8'd94, 8'd151, 8'd152, 8'd107, 8'd100, 8'd84, 8'd121, 8'd133, 8'd93, 8'd95, 8'd115, 8'd100, 8'd122, 8'd99})
) cell_0_25 (
    .clk(clk),
    .input_index(index_0_24_25),
    .input_value(value_0_24_25),
    .input_result(result_0_24_25),
    .input_enable(enable_0_24_25),
    .output_index(index_0_25_26),
    .output_value(value_0_25_26),
    .output_result(result_0_25_26),
    .output_enable(enable_0_25_26)
);

wire [10-1:0] index_0_26_27;
wire [`DATA_WIDTH-1:0] value_0_26_27;
wire [`DATA_WIDTH*4:0] result_0_26_27;
wire enable_0_26_27;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd168, 8'd164, 8'd139, 8'd169, 8'd148, 8'd83, 8'd87, 8'd132, 8'd120, 8'd136, 8'd188, 8'd159, 8'd176, 8'd141, 8'd115, 8'd161, 8'd131, 8'd95, 8'd89, 8'd169, 8'd139, 8'd85, 8'd159, 8'd119, 8'd103, 8'd118, 8'd100, 8'd83, 8'd132, 8'd154, 8'd162, 8'd113, 8'd114, 8'd167, 8'd113, 8'd74, 8'd137, 8'd89, 8'd131, 8'd67, 8'd95, 8'd123, 8'd72, 8'd104, 8'd97, 8'd120, 8'd56, 8'd73, 8'd111, 8'd57, 8'd87, 8'd75, 8'd89, 8'd127, 8'd144, 8'd115, 8'd162, 8'd81, 8'd173, 8'd125, 8'd72, 8'd129, 8'd100, 8'd81, 8'd121, 8'd123, 8'd74, 8'd64, 8'd103, 8'd108, 8'd110, 8'd73, 8'd81, 8'd128, 8'd127, 8'd93, 8'd121, 8'd114, 8'd146, 8'd124, 8'd139, 8'd80, 8'd115, 8'd146, 8'd133, 8'd165, 8'd173, 8'd125, 8'd151, 8'd118, 8'd93, 8'd102, 8'd123, 8'd106, 8'd153, 8'd95, 8'd91, 8'd140, 8'd116, 8'd134, 8'd112, 8'd122, 8'd62, 8'd58, 8'd107, 8'd149, 8'd140, 8'd66, 8'd61, 8'd118, 8'd106, 8'd97, 8'd153, 8'd171, 8'd126, 8'd142, 8'd143, 8'd87, 8'd79, 8'd142, 8'd133, 8'd167, 8'd78, 8'd133, 8'd149, 8'd90, 8'd119, 8'd94, 8'd77, 8'd155, 8'd108, 8'd86, 8'd80, 8'd142, 8'd131, 8'd157, 8'd128, 8'd119, 8'd115, 8'd72, 8'd117, 8'd144, 8'd87, 8'd163, 8'd165, 8'd116, 8'd109, 8'd160, 8'd139, 8'd149, 8'd158, 8'd106, 8'd156, 8'd61, 8'd70, 8'd90, 8'd83, 8'd152, 8'd174, 8'd127, 8'd89, 8'd155, 8'd118, 8'd143, 8'd132, 8'd114, 8'd167, 8'd115, 8'd86, 8'd103, 8'd185, 8'd157, 8'd132, 8'd127, 8'd167, 8'd169, 8'd148, 8'd148, 8'd99, 8'd105, 8'd142, 8'd137, 8'd157, 8'd135, 8'd174, 8'd99, 8'd123, 8'd183, 8'd108, 8'd74, 8'd132, 8'd177, 8'd90, 8'd110, 8'd104, 8'd130, 8'd80, 8'd119, 8'd93, 8'd140, 8'd116, 8'd131, 8'd73, 8'd147, 8'd117, 8'd104, 8'd90, 8'd90, 8'd83, 8'd101, 8'd118, 8'd172, 8'd189, 8'd142, 8'd114, 8'd176, 8'd157, 8'd146, 8'd124, 8'd101, 8'd105, 8'd168, 8'd129, 8'd131, 8'd124, 8'd158, 8'd126, 8'd98, 8'd162, 8'd74, 8'd104, 8'd92, 8'd91, 8'd68, 8'd85, 8'd80, 8'd112, 8'd99, 8'd137, 8'd135, 8'd122, 8'd144, 8'd186, 8'd170, 8'd157, 8'd161, 8'd155, 8'd81, 8'd98, 8'd167, 8'd156, 8'd112, 8'd114, 8'd160, 8'd174, 8'd198, 8'd98, 8'd98, 8'd98, 8'd101, 8'd84, 8'd88, 8'd74, 8'd69, 8'd158, 8'd103, 8'd135, 8'd135, 8'd140, 8'd93, 8'd176, 8'd168, 8'd175, 8'd154, 8'd146, 8'd156, 8'd116, 8'd107, 8'd93, 8'd148, 8'd117, 8'd209, 8'd159, 8'd163, 8'd172, 8'd164, 8'd123, 8'd105, 8'd96, 8'd118, 8'd63, 8'd76, 8'd109, 8'd120, 8'd130, 8'd130, 8'd141, 8'd163, 8'd154, 8'd72, 8'd170, 8'd161, 8'd111, 8'd150, 8'd102, 8'd95, 8'd149, 8'd88, 8'd107, 8'd171, 8'd113, 8'd136, 8'd176, 8'd158, 8'd130, 8'd150, 8'd87, 8'd128, 8'd81, 8'd82, 8'd147, 8'd136, 8'd144, 8'd91, 8'd95, 8'd133, 8'd102, 8'd110, 8'd119, 8'd87, 8'd157, 8'd136, 8'd121, 8'd83, 8'd87, 8'd124, 8'd135, 8'd135, 8'd183, 8'd183, 8'd136, 8'd165, 8'd165, 8'd143, 8'd167, 8'd84, 8'd134, 8'd71, 8'd75, 8'd147, 8'd135, 8'd88, 8'd83, 8'd85, 8'd130, 8'd153, 8'd111, 8'd100, 8'd147, 8'd83, 8'd140, 8'd157, 8'd116, 8'd83, 8'd106, 8'd203, 8'd147, 8'd183, 8'd84, 8'd109, 8'd77, 8'd94, 8'd114, 8'd95, 8'd83, 8'd125, 8'd92, 8'd106, 8'd101, 8'd57, 8'd61, 8'd93, 8'd157, 8'd87, 8'd106, 8'd157, 8'd119, 8'd157, 8'd98, 8'd156, 8'd141, 8'd139, 8'd112, 8'd128, 8'd191, 8'd172, 8'd60, 8'd135, 8'd64, 8'd95, 8'd77, 8'd56, 8'd48, 8'd51, 8'd78, 8'd113, 8'd88, 8'd118, 8'd84, 8'd104, 8'd120, 8'd72, 8'd96, 8'd98, 8'd139, 8'd137, 8'd121, 8'd140, 8'd99, 8'd133, 8'd103, 8'd157, 8'd149, 8'd121, 8'd135, 8'd61, 8'd63, 8'd104, 8'd103, 8'd81, 8'd69, 8'd83, 8'd94, 8'd74, 8'd50, 8'd150, 8'd149, 8'd119, 8'd96, 8'd70, 8'd105, 8'd109, 8'd56, 8'd128, 8'd122, 8'd166, 8'd145, 8'd146, 8'd82, 8'd179, 8'd197, 8'd129, 8'd61, 8'd149, 8'd103, 8'd120, 8'd146, 8'd68, 8'd129, 8'd165, 8'd116, 8'd82, 8'd117, 8'd130, 8'd57, 8'd95, 8'd95, 8'd136, 8'd71, 8'd92, 8'd113, 8'd169, 8'd145, 8'd152, 8'd121, 8'd78, 8'd84, 8'd173, 8'd173, 8'd97, 8'd168, 8'd114, 8'd72, 8'd98, 8'd95, 8'd123, 8'd111, 8'd91, 8'd133, 8'd152, 8'd130, 8'd107, 8'd148, 8'd140, 8'd85, 8'd162, 8'd100, 8'd100, 8'd103, 8'd173, 8'd121, 8'd108, 8'd107, 8'd177, 8'd134, 8'd181, 8'd185, 8'd135, 8'd110, 8'd97, 8'd157, 8'd88, 8'd118, 8'd171, 8'd164, 8'd113, 8'd151, 8'd125, 8'd115, 8'd96, 8'd88, 8'd126, 8'd159, 8'd84, 8'd120, 8'd71, 8'd79, 8'd178, 8'd175, 8'd182, 8'd149, 8'd122, 8'd115, 8'd134, 8'd178, 8'd135, 8'd146, 8'd91, 8'd107, 8'd91, 8'd125, 8'd134, 8'd86, 8'd124, 8'd53, 8'd127, 8'd129, 8'd100, 8'd111, 8'd130, 8'd137, 8'd93, 8'd154, 8'd165, 8'd113, 8'd153, 8'd102, 8'd153, 8'd127, 8'd88, 8'd167, 8'd99, 8'd96, 8'd157, 8'd166, 8'd129, 8'd117, 8'd137, 8'd142, 8'd90, 8'd81, 8'd63, 8'd83, 8'd107, 8'd69, 8'd137, 8'd110, 8'd61, 8'd158, 8'd113, 8'd160, 8'd140, 8'd122, 8'd173, 8'd187, 8'd170, 8'd143, 8'd114, 8'd118, 8'd110, 8'd151, 8'd102, 8'd119, 8'd156, 8'd146, 8'd90, 8'd83, 8'd86, 8'd72, 8'd74, 8'd110, 8'd94, 8'd112, 8'd72, 8'd80, 8'd111, 8'd83, 8'd107, 8'd165, 8'd163, 8'd134, 8'd111, 8'd146, 8'd137, 8'd127, 8'd163, 8'd99, 8'd82, 8'd83, 8'd121, 8'd176, 8'd204, 8'd168, 8'd139, 8'd142, 8'd144, 8'd124, 8'd142, 8'd96, 8'd108, 8'd156, 8'd149, 8'd116, 8'd91, 8'd87, 8'd152, 8'd142, 8'd164, 8'd108, 8'd74, 8'd100, 8'd154, 8'd135, 8'd163, 8'd105, 8'd140, 8'd113, 8'd131, 8'd139, 8'd163, 8'd111, 8'd133, 8'd175, 8'd178, 8'd124, 8'd108, 8'd109, 8'd106, 8'd109, 8'd133, 8'd101, 8'd92, 8'd99, 8'd64, 8'd85, 8'd120, 8'd114, 8'd90, 8'd83, 8'd90, 8'd148, 8'd83, 8'd103, 8'd125, 8'd83, 8'd140, 8'd70, 8'd71, 8'd136, 8'd152, 8'd66, 8'd103, 8'd165, 8'd129, 8'd109, 8'd128, 8'd95, 8'd86, 8'd148, 8'd91, 8'd164, 8'd108, 8'd67, 8'd94, 8'd126, 8'd88, 8'd145, 8'd163, 8'd153, 8'd136, 8'd159, 8'd144, 8'd140, 8'd129, 8'd150, 8'd111, 8'd137, 8'd113, 8'd108, 8'd103, 8'd152, 8'd122, 8'd80, 8'd144, 8'd140, 8'd102, 8'd61, 8'd72, 8'd131, 8'd71, 8'd117, 8'd112, 8'd75, 8'd147, 8'd129, 8'd103, 8'd147, 8'd102, 8'd128, 8'd83, 8'd134, 8'd145, 8'd111, 8'd88, 8'd125, 8'd138, 8'd131, 8'd120, 8'd108, 8'd129, 8'd84, 8'd108, 8'd104, 8'd127, 8'd76, 8'd124, 8'd57, 8'd71, 8'd64, 8'd126, 8'd114, 8'd97, 8'd166, 8'd126, 8'd105, 8'd99, 8'd169, 8'd132, 8'd163, 8'd127, 8'd148, 8'd122, 8'd146, 8'd107, 8'd107, 8'd95, 8'd153, 8'd126, 8'd151, 8'd124, 8'd109, 8'd98, 8'd141, 8'd94, 8'd76, 8'd109, 8'd97, 8'd71, 8'd140, 8'd156, 8'd103, 8'd169, 8'd131, 8'd109})
) cell_0_26 (
    .clk(clk),
    .input_index(index_0_25_26),
    .input_value(value_0_25_26),
    .input_result(result_0_25_26),
    .input_enable(enable_0_25_26),
    .output_index(index_0_26_27),
    .output_value(value_0_26_27),
    .output_result(result_0_26_27),
    .output_enable(enable_0_26_27)
);

wire [10-1:0] index_0_27_28;
wire [`DATA_WIDTH-1:0] value_0_27_28;
wire [`DATA_WIDTH*4:0] result_0_27_28;
wire enable_0_27_28;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd126, 8'd148, 8'd78, 8'd129, 8'd72, 8'd82, 8'd73, 8'd135, 8'd100, 8'd91, 8'd70, 8'd83, 8'd103, 8'd163, 8'd116, 8'd80, 8'd69, 8'd123, 8'd114, 8'd92, 8'd90, 8'd148, 8'd97, 8'd118, 8'd164, 8'd116, 8'd75, 8'd146, 8'd117, 8'd166, 8'd145, 8'd119, 8'd134, 8'd131, 8'd107, 8'd158, 8'd136, 8'd70, 8'd113, 8'd140, 8'd90, 8'd93, 8'd70, 8'd64, 8'd63, 8'd66, 8'd64, 8'd162, 8'd84, 8'd139, 8'd74, 8'd142, 8'd115, 8'd112, 8'd114, 8'd146, 8'd73, 8'd106, 8'd121, 8'd90, 8'd125, 8'd74, 8'd69, 8'd106, 8'd76, 8'd79, 8'd85, 8'd51, 8'd146, 8'd69, 8'd124, 8'd145, 8'd115, 8'd114, 8'd52, 8'd95, 8'd38, 8'd110, 8'd80, 8'd139, 8'd76, 8'd137, 8'd102, 8'd120, 8'd164, 8'd127, 8'd100, 8'd120, 8'd93, 8'd145, 8'd127, 8'd118, 8'd92, 8'd110, 8'd77, 8'd91, 8'd104, 8'd81, 8'd126, 8'd97, 8'd82, 8'd129, 8'd129, 8'd124, 8'd118, 8'd75, 8'd54, 8'd112, 8'd133, 8'd127, 8'd143, 8'd98, 8'd92, 8'd81, 8'd113, 8'd85, 8'd121, 8'd87, 8'd91, 8'd137, 8'd130, 8'd149, 8'd121, 8'd89, 8'd97, 8'd103, 8'd148, 8'd147, 8'd168, 8'd78, 8'd95, 8'd150, 8'd125, 8'd101, 8'd155, 8'd77, 8'd75, 8'd153, 8'd160, 8'd135, 8'd145, 8'd144, 8'd129, 8'd161, 8'd166, 8'd93, 8'd80, 8'd130, 8'd166, 8'd90, 8'd123, 8'd126, 8'd141, 8'd114, 8'd100, 8'd168, 8'd91, 8'd91, 8'd114, 8'd136, 8'd126, 8'd139, 8'd104, 8'd141, 8'd150, 8'd101, 8'd135, 8'd92, 8'd82, 8'd171, 8'd140, 8'd144, 8'd170, 8'd160, 8'd175, 8'd101, 8'd133, 8'd183, 8'd107, 8'd110, 8'd144, 8'd169, 8'd137, 8'd130, 8'd151, 8'd154, 8'd125, 8'd148, 8'd166, 8'd164, 8'd88, 8'd159, 8'd105, 8'd129, 8'd132, 8'd165, 8'd135, 8'd152, 8'd104, 8'd117, 8'd109, 8'd182, 8'd157, 8'd87, 8'd118, 8'd142, 8'd115, 8'd147, 8'd168, 8'd104, 8'd162, 8'd99, 8'd168, 8'd122, 8'd107, 8'd153, 8'd185, 8'd119, 8'd133, 8'd124, 8'd85, 8'd165, 8'd158, 8'd93, 8'd139, 8'd105, 8'd144, 8'd170, 8'd111, 8'd123, 8'd158, 8'd112, 8'd126, 8'd132, 8'd78, 8'd173, 8'd169, 8'd160, 8'd118, 8'd158, 8'd141, 8'd156, 8'd120, 8'd183, 8'd146, 8'd115, 8'd81, 8'd133, 8'd129, 8'd77, 8'd90, 8'd94, 8'd100, 8'd102, 8'd172, 8'd188, 8'd147, 8'd137, 8'd127, 8'd118, 8'd112, 8'd136, 8'd118, 8'd75, 8'd126, 8'd76, 8'd112, 8'd164, 8'd162, 8'd180, 8'd114, 8'd120, 8'd136, 8'd126, 8'd78, 8'd153, 8'd95, 8'd142, 8'd86, 8'd133, 8'd174, 8'd145, 8'd159, 8'd117, 8'd174, 8'd171, 8'd139, 8'd130, 8'd63, 8'd130, 8'd109, 8'd105, 8'd63, 8'd154, 8'd139, 8'd104, 8'd156, 8'd150, 8'd124, 8'd97, 8'd143, 8'd129, 8'd134, 8'd142, 8'd146, 8'd111, 8'd95, 8'd144, 8'd175, 8'd193, 8'd179, 8'd136, 8'd166, 8'd108, 8'd158, 8'd108, 8'd58, 8'd69, 8'd90, 8'd75, 8'd123, 8'd108, 8'd152, 8'd159, 8'd135, 8'd77, 8'd75, 8'd111, 8'd112, 8'd102, 8'd130, 8'd137, 8'd91, 8'd117, 8'd161, 8'd150, 8'd184, 8'd110, 8'd137, 8'd159, 8'd131, 8'd153, 8'd94, 8'd155, 8'd82, 8'd122, 8'd47, 8'd131, 8'd121, 8'd107, 8'd103, 8'd103, 8'd138, 8'd152, 8'd147, 8'd111, 8'd72, 8'd95, 8'd109, 8'd69, 8'd98, 8'd133, 8'd148, 8'd104, 8'd93, 8'd140, 8'd146, 8'd121, 8'd126, 8'd111, 8'd137, 8'd57, 8'd84, 8'd73, 8'd137, 8'd114, 8'd137, 8'd168, 8'd166, 8'd147, 8'd122, 8'd132, 8'd109, 8'd130, 8'd80, 8'd91, 8'd103, 8'd106, 8'd72, 8'd169, 8'd132, 8'd145, 8'd157, 8'd105, 8'd101, 8'd169, 8'd146, 8'd81, 8'd70, 8'd120, 8'd127, 8'd64, 8'd93, 8'd96, 8'd128, 8'd139, 8'd102, 8'd127, 8'd139, 8'd72, 8'd61, 8'd53, 8'd73, 8'd105, 8'd58, 8'd79, 8'd105, 8'd127, 8'd84, 8'd111, 8'd131, 8'd124, 8'd103, 8'd216, 8'd130, 8'd123, 8'd126, 8'd111, 8'd164, 8'd130, 8'd108, 8'd91, 8'd165, 8'd145, 8'd112, 8'd100, 8'd59, 8'd68, 8'd98, 8'd80, 8'd64, 8'd105, 8'd92, 8'd76, 8'd118, 8'd108, 8'd165, 8'd117, 8'd132, 8'd75, 8'd135, 8'd91, 8'd188, 8'd104, 8'd146, 8'd100, 8'd157, 8'd123, 8'd126, 8'd131, 8'd98, 8'd131, 8'd70, 8'd90, 8'd51, 8'd91, 8'd53, 8'd56, 8'd87, 8'd146, 8'd67, 8'd146, 8'd166, 8'd178, 8'd95, 8'd120, 8'd151, 8'd114, 8'd38, 8'd53, 8'd105, 8'd105, 8'd154, 8'd172, 8'd111, 8'd99, 8'd145, 8'd101, 8'd127, 8'd169, 8'd168, 8'd128, 8'd124, 8'd119, 8'd93, 8'd143, 8'd111, 8'd167, 8'd110, 8'd165, 8'd151, 8'd136, 8'd136, 8'd117, 8'd120, 8'd103, 8'd124, 8'd127, 8'd117, 8'd71, 8'd131, 8'd105, 8'd99, 8'd72, 8'd146, 8'd143, 8'd130, 8'd122, 8'd131, 8'd146, 8'd129, 8'd114, 8'd67, 8'd85, 8'd162, 8'd133, 8'd103, 8'd109, 8'd103, 8'd81, 8'd80, 8'd85, 8'd166, 8'd162, 8'd53, 8'd64, 8'd74, 8'd131, 8'd70, 8'd95, 8'd128, 8'd119, 8'd104, 8'd174, 8'd186, 8'd162, 8'd154, 8'd73, 8'd107, 8'd126, 8'd78, 8'd94, 8'd128, 8'd115, 8'd170, 8'd177, 8'd120, 8'd63, 8'd142, 8'd100, 8'd94, 8'd160, 8'd55, 8'd107, 8'd88, 8'd160, 8'd82, 8'd157, 8'd115, 8'd73, 8'd122, 8'd141, 8'd111, 8'd77, 8'd141, 8'd95, 8'd96, 8'd125, 8'd154, 8'd79, 8'd154, 8'd118, 8'd140, 8'd114, 8'd85, 8'd101, 8'd132, 8'd133, 8'd77, 8'd62, 8'd96, 8'd46, 8'd129, 8'd143, 8'd117, 8'd139, 8'd142, 8'd111, 8'd99, 8'd136, 8'd129, 8'd100, 8'd79, 8'd150, 8'd165, 8'd117, 8'd114, 8'd109, 8'd128, 8'd92, 8'd143, 8'd116, 8'd112, 8'd81, 8'd128, 8'd161, 8'd108, 8'd64, 8'd72, 8'd139, 8'd90, 8'd97, 8'd123, 8'd76, 8'd82, 8'd104, 8'd87, 8'd137, 8'd122, 8'd112, 8'd124, 8'd148, 8'd143, 8'd97, 8'd146, 8'd157, 8'd151, 8'd131, 8'd174, 8'd102, 8'd117, 8'd128, 8'd87, 8'd110, 8'd95, 8'd118, 8'd91, 8'd125, 8'd122, 8'd114, 8'd70, 8'd105, 8'd161, 8'd123, 8'd154, 8'd122, 8'd133, 8'd146, 8'd184, 8'd170, 8'd115, 8'd191, 8'd146, 8'd196, 8'd119, 8'd165, 8'd99, 8'd154, 8'd178, 8'd93, 8'd165, 8'd123, 8'd119, 8'd147, 8'd73, 8'd166, 8'd160, 8'd76, 8'd103, 8'd100, 8'd150, 8'd122, 8'd113, 8'd188, 8'd108, 8'd170, 8'd155, 8'd197, 8'd175, 8'd202, 8'd134, 8'd111, 8'd114, 8'd119, 8'd101, 8'd153, 8'd101, 8'd105, 8'd158, 8'd144, 8'd103, 8'd115, 8'd138, 8'd123, 8'd115, 8'd108, 8'd87, 8'd136, 8'd164, 8'd122, 8'd115, 8'd132, 8'd218, 8'd196, 8'd168, 8'd211, 8'd155, 8'd137, 8'd118, 8'd136, 8'd100, 8'd108, 8'd101, 8'd162, 8'd88, 8'd134, 8'd166, 8'd164, 8'd77, 8'd76, 8'd148, 8'd79, 8'd162, 8'd178, 8'd178, 8'd150, 8'd121, 8'd97, 8'd131, 8'd192, 8'd115, 8'd141, 8'd194, 8'd155, 8'd124, 8'd125, 8'd172, 8'd107, 8'd97, 8'd148, 8'd137, 8'd113, 8'd110, 8'd106, 8'd134, 8'd135, 8'd119, 8'd92, 8'd163, 8'd132, 8'd149, 8'd103, 8'd106, 8'd119, 8'd94, 8'd79, 8'd141, 8'd162, 8'd149, 8'd145, 8'd123, 8'd84, 8'd121, 8'd165, 8'd95, 8'd84, 8'd159, 8'd77, 8'd100, 8'd100, 8'd137, 8'd104, 8'd78, 8'd167})
) cell_0_27 (
    .clk(clk),
    .input_index(index_0_26_27),
    .input_value(value_0_26_27),
    .input_result(result_0_26_27),
    .input_enable(enable_0_26_27),
    .output_index(index_0_27_28),
    .output_value(value_0_27_28),
    .output_result(result_0_27_28),
    .output_enable(enable_0_27_28)
);

wire [10-1:0] index_0_28_29;
wire [`DATA_WIDTH-1:0] value_0_28_29;
wire [`DATA_WIDTH*4:0] result_0_28_29;
wire enable_0_28_29;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd133, 8'd166, 8'd117, 8'd105, 8'd163, 8'd162, 8'd171, 8'd165, 8'd165, 8'd104, 8'd170, 8'd126, 8'd120, 8'd146, 8'd158, 8'd169, 8'd162, 8'd190, 8'd115, 8'd92, 8'd143, 8'd158, 8'd131, 8'd118, 8'd162, 8'd161, 8'd82, 8'd88, 8'd106, 8'd123, 8'd148, 8'd155, 8'd115, 8'd126, 8'd97, 8'd145, 8'd127, 8'd154, 8'd164, 8'd134, 8'd169, 8'd137, 8'd157, 8'd131, 8'd210, 8'd155, 8'd121, 8'd201, 8'd190, 8'd169, 8'd141, 8'd128, 8'd151, 8'd144, 8'd168, 8'd149, 8'd164, 8'd158, 8'd165, 8'd159, 8'd99, 8'd95, 8'd164, 8'd195, 8'd135, 8'd193, 8'd200, 8'd187, 8'd154, 8'd158, 8'd121, 8'd160, 8'd157, 8'd191, 8'd221, 8'd161, 8'd179, 8'd204, 8'd196, 8'd108, 8'd146, 8'd84, 8'd159, 8'd148, 8'd169, 8'd111, 8'd61, 8'd119, 8'd109, 8'd70, 8'd115, 8'd137, 8'd62, 8'd162, 8'd94, 8'd95, 8'd110, 8'd64, 8'd124, 8'd160, 8'd109, 8'd118, 8'd100, 8'd201, 8'd193, 8'd213, 8'd194, 8'd130, 8'd187, 8'd124, 8'd70, 8'd95, 8'd121, 8'd113, 8'd144, 8'd88, 8'd125, 8'd53, 8'd45, 8'd47, 8'd111, 8'd97, 8'd155, 8'd95, 8'd148, 8'd68, 8'd142, 8'd94, 8'd138, 8'd117, 8'd148, 8'd155, 8'd165, 8'd145, 8'd199, 8'd108, 8'd176, 8'd81, 8'd145, 8'd150, 8'd95, 8'd116, 8'd83, 8'd91, 8'd85, 8'd115, 8'd97, 8'd111, 8'd91, 8'd155, 8'd115, 8'd143, 8'd136, 8'd76, 8'd80, 8'd124, 8'd153, 8'd120, 8'd116, 8'd95, 8'd87, 8'd148, 8'd182, 8'd84, 8'd112, 8'd142, 8'd115, 8'd80, 8'd161, 8'd109, 8'd145, 8'd159, 8'd69, 8'd111, 8'd87, 8'd153, 8'd62, 8'd165, 8'd150, 8'd151, 8'd79, 8'd169, 8'd100, 8'd123, 8'd140, 8'd156, 8'd148, 8'd91, 8'd110, 8'd170, 8'd97, 8'd127, 8'd164, 8'd131, 8'd166, 8'd167, 8'd148, 8'd101, 8'd95, 8'd111, 8'd68, 8'd132, 8'd68, 8'd101, 8'd114, 8'd148, 8'd79, 8'd138, 8'd165, 8'd134, 8'd170, 8'd123, 8'd86, 8'd175, 8'd107, 8'd76, 8'd150, 8'd163, 8'd139, 8'd145, 8'd95, 8'd107, 8'd110, 8'd102, 8'd90, 8'd64, 8'd111, 8'd155, 8'd88, 8'd77, 8'd84, 8'd78, 8'd124, 8'd134, 8'd154, 8'd133, 8'd143, 8'd159, 8'd168, 8'd155, 8'd103, 8'd93, 8'd67, 8'd63, 8'd135, 8'd122, 8'd113, 8'd110, 8'd178, 8'd99, 8'd108, 8'd167, 8'd111, 8'd140, 8'd96, 8'd92, 8'd133, 8'd88, 8'd149, 8'd134, 8'd143, 8'd90, 8'd135, 8'd95, 8'd151, 8'd71, 8'd106, 8'd57, 8'd63, 8'd136, 8'd78, 8'd62, 8'd66, 8'd106, 8'd169, 8'd107, 8'd185, 8'd152, 8'd164, 8'd132, 8'd99, 8'd141, 8'd92, 8'd76, 8'd129, 8'd131, 8'd134, 8'd171, 8'd128, 8'd105, 8'd82, 8'd121, 8'd87, 8'd156, 8'd128, 8'd106, 8'd103, 8'd74, 8'd66, 8'd60, 8'd77, 8'd161, 8'd117, 8'd99, 8'd124, 8'd176, 8'd179, 8'd148, 8'd66, 8'd100, 8'd62, 8'd115, 8'd92, 8'd97, 8'd92, 8'd184, 8'd134, 8'd164, 8'd77, 8'd64, 8'd100, 8'd138, 8'd130, 8'd70, 8'd150, 8'd58, 8'd72, 8'd70, 8'd126, 8'd111, 8'd146, 8'd132, 8'd140, 8'd98, 8'd125, 8'd151, 8'd98, 8'd48, 8'd120, 8'd154, 8'd92, 8'd105, 8'd102, 8'd111, 8'd143, 8'd88, 8'd77, 8'd78, 8'd81, 8'd118, 8'd110, 8'd79, 8'd130, 8'd113, 8'd104, 8'd89, 8'd122, 8'd71, 8'd77, 8'd91, 8'd82, 8'd175, 8'd166, 8'd115, 8'd133, 8'd81, 8'd75, 8'd162, 8'd132, 8'd118, 8'd135, 8'd95, 8'd114, 8'd124, 8'd97, 8'd101, 8'd126, 8'd108, 8'd133, 8'd34, 8'd105, 8'd56, 8'd131, 8'd68, 8'd146, 8'd69, 8'd79, 8'd75, 8'd157, 8'd95, 8'd99, 8'd155, 8'd152, 8'd120, 8'd55, 8'd81, 8'd120, 8'd72, 8'd109, 8'd102, 8'd91, 8'd118, 8'd87, 8'd112, 8'd123, 8'd150, 8'd124, 8'd106, 8'd57, 8'd77, 8'd141, 8'd147, 8'd153, 8'd72, 8'd80, 8'd99, 8'd103, 8'd111, 8'd102, 8'd121, 8'd169, 8'd121, 8'd135, 8'd129, 8'd96, 8'd121, 8'd83, 8'd117, 8'd95, 8'd143, 8'd134, 8'd102, 8'd145, 8'd140, 8'd92, 8'd82, 8'd74, 8'd121, 8'd148, 8'd129, 8'd73, 8'd155, 8'd129, 8'd124, 8'd191, 8'd108, 8'd145, 8'd108, 8'd96, 8'd76, 8'd127, 8'd114, 8'd135, 8'd96, 8'd71, 8'd143, 8'd102, 8'd141, 8'd127, 8'd103, 8'd111, 8'd119, 8'd103, 8'd82, 8'd103, 8'd115, 8'd90, 8'd88, 8'd81, 8'd132, 8'd125, 8'd98, 8'd187, 8'd164, 8'd159, 8'd123, 8'd68, 8'd62, 8'd83, 8'd129, 8'd109, 8'd138, 8'd142, 8'd161, 8'd95, 8'd162, 8'd175, 8'd192, 8'd201, 8'd190, 8'd123, 8'd135, 8'd79, 8'd57, 8'd45, 8'd64, 8'd139, 8'd101, 8'd142, 8'd159, 8'd108, 8'd130, 8'd121, 8'd163, 8'd112, 8'd52, 8'd33, 8'd39, 8'd92, 8'd104, 8'd99, 8'd96, 8'd98, 8'd134, 8'd149, 8'd195, 8'd140, 8'd160, 8'd151, 8'd82, 8'd153, 8'd137, 8'd112, 8'd74, 8'd129, 8'd160, 8'd135, 8'd187, 8'd186, 8'd163, 8'd109, 8'd128, 8'd132, 8'd58, 8'd3, 8'd57, 8'd49, 8'd137, 8'd75, 8'd126, 8'd104, 8'd111, 8'd190, 8'd142, 8'd129, 8'd197, 8'd143, 8'd150, 8'd153, 8'd172, 8'd143, 8'd130, 8'd88, 8'd175, 8'd135, 8'd177, 8'd121, 8'd137, 8'd124, 8'd156, 8'd70, 8'd73, 8'd105, 8'd106, 8'd111, 8'd109, 8'd49, 8'd117, 8'd70, 8'd138, 8'd190, 8'd128, 8'd180, 8'd129, 8'd123, 8'd206, 8'd111, 8'd180, 8'd105, 8'd159, 8'd148, 8'd146, 8'd148, 8'd130, 8'd105, 8'd140, 8'd106, 8'd132, 8'd116, 8'd103, 8'd56, 8'd81, 8'd74, 8'd40, 8'd90, 8'd67, 8'd126, 8'd130, 8'd86, 8'd116, 8'd179, 8'd191, 8'd166, 8'd127, 8'd158, 8'd152, 8'd133, 8'd111, 8'd105, 8'd85, 8'd109, 8'd175, 8'd169, 8'd127, 8'd78, 8'd165, 8'd120, 8'd78, 8'd95, 8'd94, 8'd60, 8'd106, 8'd54, 8'd117, 8'd107, 8'd131, 8'd102, 8'd45, 8'd76, 8'd149, 8'd111, 8'd132, 8'd101, 8'd74, 8'd88, 8'd125, 8'd82, 8'd110, 8'd121, 8'd153, 8'd105, 8'd104, 8'd133, 8'd146, 8'd140, 8'd171, 8'd134, 8'd88, 8'd139, 8'd94, 8'd85, 8'd88, 8'd141, 8'd119, 8'd158, 8'd133, 8'd92, 8'd100, 8'd112, 8'd112, 8'd147, 8'd90, 8'd127, 8'd140, 8'd80, 8'd118, 8'd109, 8'd91, 8'd110, 8'd164, 8'd82, 8'd97, 8'd117, 8'd81, 8'd162, 8'd116, 8'd124, 8'd165, 8'd162, 8'd151, 8'd119, 8'd128, 8'd106, 8'd155, 8'd196, 8'd146, 8'd190, 8'd160, 8'd173, 8'd163, 8'd105, 8'd186, 8'd175, 8'd118, 8'd146, 8'd75, 8'd162, 8'd82, 8'd153, 8'd128, 8'd88, 8'd122, 8'd160, 8'd98, 8'd101, 8'd181, 8'd143, 8'd156, 8'd117, 8'd96, 8'd154, 8'd155, 8'd178, 8'd169, 8'd122, 8'd196, 8'd165, 8'd189, 8'd193, 8'd192, 8'd118, 8'd124, 8'd108, 8'd114, 8'd84, 8'd95, 8'd151, 8'd89, 8'd76, 8'd106, 8'd88, 8'd169, 8'd93, 8'd147, 8'd157, 8'd149, 8'd92, 8'd179, 8'd138, 8'd148, 8'd191, 8'd103, 8'd143, 8'd136, 8'd139, 8'd107, 8'd162, 8'd125, 8'd147, 8'd132, 8'd120, 8'd82, 8'd124, 8'd111, 8'd80, 8'd106, 8'd116, 8'd156, 8'd104, 8'd89, 8'd117, 8'd81, 8'd102, 8'd167, 8'd166, 8'd109, 8'd151, 8'd166, 8'd92, 8'd104, 8'd116, 8'd110, 8'd136, 8'd129, 8'd152, 8'd100, 8'd97, 8'd141, 8'd88, 8'd91, 8'd120, 8'd81, 8'd125, 8'd155})
) cell_0_28 (
    .clk(clk),
    .input_index(index_0_27_28),
    .input_value(value_0_27_28),
    .input_result(result_0_27_28),
    .input_enable(enable_0_27_28),
    .output_index(index_0_28_29),
    .output_value(value_0_28_29),
    .output_result(result_0_28_29),
    .output_enable(enable_0_28_29)
);

wire [10-1:0] index_0_29_30;
wire [`DATA_WIDTH-1:0] value_0_29_30;
wire [`DATA_WIDTH*4:0] result_0_29_30;
wire enable_0_29_30;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd90, 8'd134, 8'd138, 8'd151, 8'd125, 8'd147, 8'd112, 8'd89, 8'd108, 8'd76, 8'd135, 8'd168, 8'd94, 8'd155, 8'd103, 8'd153, 8'd101, 8'd126, 8'd98, 8'd97, 8'd138, 8'd168, 8'd158, 8'd137, 8'd107, 8'd131, 8'd87, 8'd144, 8'd160, 8'd130, 8'd146, 8'd162, 8'd85, 8'd113, 8'd93, 8'd119, 8'd79, 8'd87, 8'd72, 8'd134, 8'd111, 8'd49, 8'd72, 8'd83, 8'd118, 8'd122, 8'd64, 8'd107, 8'd89, 8'd121, 8'd100, 8'd98, 8'd77, 8'd84, 8'd165, 8'd153, 8'd130, 8'd166, 8'd101, 8'd111, 8'd162, 8'd125, 8'd50, 8'd97, 8'd60, 8'd58, 8'd65, 8'd150, 8'd145, 8'd124, 8'd120, 8'd88, 8'd90, 8'd106, 8'd103, 8'd130, 8'd128, 8'd69, 8'd110, 8'd121, 8'd140, 8'd153, 8'd163, 8'd164, 8'd141, 8'd174, 8'd79, 8'd67, 8'd135, 8'd131, 8'd152, 8'd160, 8'd162, 8'd101, 8'd100, 8'd138, 8'd161, 8'd143, 8'd141, 8'd154, 8'd152, 8'd133, 8'd109, 8'd78, 8'd123, 8'd140, 8'd165, 8'd108, 8'd181, 8'd89, 8'd159, 8'd152, 8'd129, 8'd166, 8'd146, 8'd104, 8'd86, 8'd143, 8'd160, 8'd82, 8'd109, 8'd132, 8'd156, 8'd155, 8'd171, 8'd139, 8'd110, 8'd138, 8'd116, 8'd149, 8'd103, 8'd87, 8'd136, 8'd99, 8'd109, 8'd193, 8'd94, 8'd90, 8'd76, 8'd95, 8'd160, 8'd147, 8'd140, 8'd90, 8'd123, 8'd113, 8'd155, 8'd162, 8'd157, 8'd145, 8'd118, 8'd159, 8'd105, 8'd124, 8'd118, 8'd86, 8'd136, 8'd131, 8'd123, 8'd121, 8'd116, 8'd147, 8'd139, 8'd179, 8'd92, 8'd125, 8'd143, 8'd82, 8'd149, 8'd127, 8'd137, 8'd143, 8'd101, 8'd105, 8'd114, 8'd92, 8'd167, 8'd152, 8'd175, 8'd124, 8'd89, 8'd105, 8'd137, 8'd78, 8'd104, 8'd91, 8'd88, 8'd133, 8'd70, 8'd115, 8'd64, 8'd175, 8'd136, 8'd82, 8'd81, 8'd151, 8'd84, 8'd108, 8'd100, 8'd71, 8'd73, 8'd113, 8'd163, 8'd100, 8'd92, 8'd150, 8'd124, 8'd173, 8'd119, 8'd127, 8'd108, 8'd116, 8'd128, 8'd91, 8'd117, 8'd76, 8'd95, 8'd83, 8'd154, 8'd80, 8'd102, 8'd96, 8'd96, 8'd108, 8'd81, 8'd122, 8'd136, 8'd121, 8'd105, 8'd109, 8'd164, 8'd71, 8'd124, 8'd166, 8'd79, 8'd118, 8'd148, 8'd153, 8'd123, 8'd143, 8'd143, 8'd110, 8'd134, 8'd79, 8'd102, 8'd116, 8'd100, 8'd106, 8'd92, 8'd175, 8'd91, 8'd125, 8'd72, 8'd130, 8'd49, 8'd81, 8'd92, 8'd123, 8'd89, 8'd77, 8'd126, 8'd154, 8'd93, 8'd94, 8'd177, 8'd113, 8'd127, 8'd137, 8'd108, 8'd97, 8'd111, 8'd64, 8'd146, 8'd83, 8'd119, 8'd165, 8'd82, 8'd150, 8'd147, 8'd125, 8'd142, 8'd140, 8'd112, 8'd130, 8'd105, 8'd92, 8'd96, 8'd162, 8'd104, 8'd124, 8'd166, 8'd107, 8'd96, 8'd180, 8'd135, 8'd106, 8'd107, 8'd132, 8'd75, 8'd120, 8'd163, 8'd95, 8'd107, 8'd83, 8'd78, 8'd116, 8'd86, 8'd96, 8'd134, 8'd75, 8'd97, 8'd144, 8'd169, 8'd157, 8'd162, 8'd139, 8'd139, 8'd116, 8'd165, 8'd168, 8'd112, 8'd112, 8'd101, 8'd126, 8'd107, 8'd113, 8'd106, 8'd144, 8'd163, 8'd74, 8'd95, 8'd57, 8'd151, 8'd99, 8'd172, 8'd103, 8'd89, 8'd128, 8'd130, 8'd144, 8'd112, 8'd87, 8'd152, 8'd124, 8'd84, 8'd120, 8'd147, 8'd130, 8'd87, 8'd158, 8'd108, 8'd103, 8'd163, 8'd109, 8'd145, 8'd162, 8'd80, 8'd119, 8'd112, 8'd98, 8'd155, 8'd96, 8'd165, 8'd161, 8'd104, 8'd132, 8'd141, 8'd112, 8'd119, 8'd100, 8'd134, 8'd113, 8'd80, 8'd104, 8'd162, 8'd168, 8'd154, 8'd113, 8'd157, 8'd141, 8'd175, 8'd117, 8'd89, 8'd141, 8'd169, 8'd82, 8'd120, 8'd93, 8'd144, 8'd95, 8'd96, 8'd88, 8'd86, 8'd165, 8'd152, 8'd138, 8'd130, 8'd62, 8'd145, 8'd109, 8'd113, 8'd157, 8'd119, 8'd147, 8'd96, 8'd79, 8'd154, 8'd99, 8'd192, 8'd101, 8'd119, 8'd161, 8'd99, 8'd106, 8'd124, 8'd115, 8'd83, 8'd108, 8'd139, 8'd159, 8'd139, 8'd135, 8'd143, 8'd127, 8'd68, 8'd59, 8'd109, 8'd90, 8'd61, 8'd132, 8'd69, 8'd72, 8'd120, 8'd64, 8'd118, 8'd188, 8'd116, 8'd142, 8'd133, 8'd162, 8'd162, 8'd101, 8'd139, 8'd156, 8'd108, 8'd144, 8'd99, 8'd138, 8'd143, 8'd116, 8'd134, 8'd88, 8'd133, 8'd54, 8'd76, 8'd84, 8'd93, 8'd75, 8'd138, 8'd164, 8'd91, 8'd63, 8'd134, 8'd140, 8'd147, 8'd138, 8'd116, 8'd93, 8'd124, 8'd104, 8'd94, 8'd74, 8'd139, 8'd134, 8'd141, 8'd109, 8'd137, 8'd184, 8'd180, 8'd168, 8'd84, 8'd89, 8'd116, 8'd64, 8'd112, 8'd146, 8'd157, 8'd107, 8'd65, 8'd111, 8'd108, 8'd133, 8'd116, 8'd84, 8'd98, 8'd174, 8'd120, 8'd105, 8'd99, 8'd94, 8'd152, 8'd152, 8'd156, 8'd117, 8'd151, 8'd187, 8'd132, 8'd144, 8'd166, 8'd109, 8'd171, 8'd147, 8'd165, 8'd122, 8'd91, 8'd96, 8'd116, 8'd62, 8'd104, 8'd96, 8'd89, 8'd103, 8'd118, 8'd158, 8'd167, 8'd142, 8'd78, 8'd119, 8'd167, 8'd183, 8'd85, 8'd101, 8'd148, 8'd154, 8'd140, 8'd182, 8'd168, 8'd121, 8'd157, 8'd127, 8'd80, 8'd144, 8'd92, 8'd82, 8'd65, 8'd68, 8'd138, 8'd128, 8'd140, 8'd123, 8'd104, 8'd119, 8'd145, 8'd114, 8'd133, 8'd111, 8'd117, 8'd98, 8'd107, 8'd105, 8'd135, 8'd103, 8'd195, 8'd170, 8'd123, 8'd142, 8'd150, 8'd81, 8'd132, 8'd147, 8'd150, 8'd47, 8'd59, 8'd71, 8'd55, 8'd71, 8'd64, 8'd125, 8'd118, 8'd103, 8'd169, 8'd163, 8'd152, 8'd134, 8'd146, 8'd167, 8'd106, 8'd97, 8'd160, 8'd176, 8'd145, 8'd188, 8'd179, 8'd164, 8'd96, 8'd156, 8'd119, 8'd135, 8'd127, 8'd130, 8'd114, 8'd106, 8'd116, 8'd147, 8'd133, 8'd75, 8'd81, 8'd87, 8'd107, 8'd139, 8'd162, 8'd109, 8'd138, 8'd130, 8'd174, 8'd90, 8'd94, 8'd155, 8'd143, 8'd159, 8'd184, 8'd168, 8'd103, 8'd154, 8'd151, 8'd153, 8'd104, 8'd102, 8'd71, 8'd97, 8'd67, 8'd119, 8'd83, 8'd92, 8'd120, 8'd148, 8'd115, 8'd127, 8'd148, 8'd104, 8'd133, 8'd130, 8'd117, 8'd107, 8'd77, 8'd92, 8'd143, 8'd152, 8'd99, 8'd139, 8'd105, 8'd107, 8'd102, 8'd176, 8'd141, 8'd157, 8'd78, 8'd100, 8'd140, 8'd83, 8'd119, 8'd154, 8'd131, 8'd103, 8'd160, 8'd96, 8'd80, 8'd109, 8'd135, 8'd124, 8'd91, 8'd112, 8'd74, 8'd102, 8'd111, 8'd102, 8'd119, 8'd128, 8'd107, 8'd113, 8'd166, 8'd144, 8'd80, 8'd96, 8'd152, 8'd58, 8'd125, 8'd83, 8'd116, 8'd123, 8'd133, 8'd130, 8'd73, 8'd63, 8'd125, 8'd111, 8'd122, 8'd70, 8'd155, 8'd75, 8'd85, 8'd127, 8'd161, 8'd65, 8'd93, 8'd103, 8'd75, 8'd146, 8'd97, 8'd67, 8'd84, 8'd61, 8'd34, 8'd31, 8'd60, 8'd16, 8'd44, 8'd38, 8'd92, 8'd113, 8'd109, 8'd63, 8'd153, 8'd73, 8'd162, 8'd157, 8'd133, 8'd82, 8'd110, 8'd81, 8'd117, 8'd157, 8'd159, 8'd139, 8'd91, 8'd128, 8'd131, 8'd133, 8'd73, 8'd140, 8'd55, 8'd95, 8'd138, 8'd89, 8'd67, 8'd107, 8'd65, 8'd116, 8'd141, 8'd141, 8'd135, 8'd161, 8'd125, 8'd72, 8'd88, 8'd148, 8'd105, 8'd118, 8'd82, 8'd120, 8'd158, 8'd87, 8'd117, 8'd163, 8'd74, 8'd102, 8'd70, 8'd117, 8'd123, 8'd165, 8'd156, 8'd68, 8'd123, 8'd150, 8'd123, 8'd102, 8'd109, 8'd73, 8'd160, 8'd146, 8'd119, 8'd87, 8'd150, 8'd137})
) cell_0_29 (
    .clk(clk),
    .input_index(index_0_28_29),
    .input_value(value_0_28_29),
    .input_result(result_0_28_29),
    .input_enable(enable_0_28_29),
    .output_index(index_0_29_30),
    .output_value(value_0_29_30),
    .output_result(result_0_29_30),
    .output_enable(enable_0_29_30)
);

wire [10-1:0] index_0_30_31;
wire [`DATA_WIDTH-1:0] value_0_30_31;
wire [`DATA_WIDTH*4:0] result_0_30_31;
wire enable_0_30_31;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd88, 8'd106, 8'd159, 8'd140, 8'd178, 8'd131, 8'd165, 8'd92, 8'd148, 8'd126, 8'd178, 8'd107, 8'd155, 8'd164, 8'd116, 8'd177, 8'd126, 8'd167, 8'd152, 8'd168, 8'd172, 8'd170, 8'd177, 8'd169, 8'd101, 8'd141, 8'd141, 8'd122, 8'd90, 8'd74, 8'd118, 8'd113, 8'd107, 8'd133, 8'd147, 8'd119, 8'd160, 8'd137, 8'd154, 8'd167, 8'd108, 8'd115, 8'd107, 8'd153, 8'd165, 8'd90, 8'd120, 8'd89, 8'd148, 8'd109, 8'd124, 8'd153, 8'd107, 8'd145, 8'd88, 8'd79, 8'd102, 8'd141, 8'd121, 8'd136, 8'd97, 8'd81, 8'd94, 8'd145, 8'd151, 8'd85, 8'd184, 8'd173, 8'd163, 8'd128, 8'd196, 8'd197, 8'd136, 8'd171, 8'd104, 8'd174, 8'd107, 8'd177, 8'd190, 8'd191, 8'd137, 8'd102, 8'd128, 8'd78, 8'd150, 8'd97, 8'd161, 8'd164, 8'd77, 8'd77, 8'd143, 8'd75, 8'd68, 8'd70, 8'd165, 8'd82, 8'd106, 8'd160, 8'd149, 8'd91, 8'd89, 8'd155, 8'd167, 8'd173, 8'd113, 8'd193, 8'd203, 8'd110, 8'd159, 8'd76, 8'd93, 8'd142, 8'd129, 8'd111, 8'd131, 8'd160, 8'd100, 8'd148, 8'd98, 8'd103, 8'd142, 8'd100, 8'd116, 8'd89, 8'd91, 8'd61, 8'd59, 8'd69, 8'd118, 8'd119, 8'd146, 8'd127, 8'd159, 8'd128, 8'd112, 8'd185, 8'd96, 8'd100, 8'd71, 8'd111, 8'd167, 8'd132, 8'd116, 8'd122, 8'd148, 8'd125, 8'd127, 8'd102, 8'd144, 8'd151, 8'd89, 8'd117, 8'd82, 8'd93, 8'd157, 8'd75, 8'd106, 8'd130, 8'd119, 8'd169, 8'd126, 8'd151, 8'd140, 8'd138, 8'd157, 8'd102, 8'd96, 8'd138, 8'd91, 8'd102, 8'd134, 8'd109, 8'd92, 8'd160, 8'd131, 8'd95, 8'd141, 8'd152, 8'd151, 8'd144, 8'd86, 8'd114, 8'd171, 8'd171, 8'd165, 8'd146, 8'd160, 8'd141, 8'd106, 8'd120, 8'd170, 8'd153, 8'd100, 8'd111, 8'd92, 8'd113, 8'd149, 8'd151, 8'd120, 8'd98, 8'd158, 8'd98, 8'd72, 8'd164, 8'd145, 8'd137, 8'd90, 8'd149, 8'd175, 8'd177, 8'd156, 8'd186, 8'd179, 8'd102, 8'd121, 8'd165, 8'd162, 8'd84, 8'd124, 8'd148, 8'd149, 8'd91, 8'd97, 8'd71, 8'd99, 8'd188, 8'd181, 8'd169, 8'd139, 8'd153, 8'd146, 8'd104, 8'd134, 8'd169, 8'd105, 8'd79, 8'd147, 8'd139, 8'd103, 8'd119, 8'd191, 8'd96, 8'd106, 8'd172, 8'd166, 8'd132, 8'd130, 8'd163, 8'd111, 8'd123, 8'd169, 8'd148, 8'd142, 8'd194, 8'd139, 8'd121, 8'd122, 8'd127, 8'd112, 8'd109, 8'd110, 8'd111, 8'd93, 8'd140, 8'd141, 8'd130, 8'd95, 8'd106, 8'd101, 8'd164, 8'd92, 8'd94, 8'd88, 8'd147, 8'd157, 8'd178, 8'd149, 8'd132, 8'd92, 8'd167, 8'd123, 8'd161, 8'd175, 8'd161, 8'd150, 8'd133, 8'd187, 8'd97, 8'd170, 8'd134, 8'd123, 8'd71, 8'd145, 8'd77, 8'd124, 8'd130, 8'd75, 8'd71, 8'd121, 8'd88, 8'd147, 8'd139, 8'd182, 8'd191, 8'd159, 8'd113, 8'd116, 8'd124, 8'd87, 8'd185, 8'd216, 8'd180, 8'd140, 8'd109, 8'd190, 8'd185, 8'd166, 8'd145, 8'd129, 8'd143, 8'd137, 8'd124, 8'd91, 8'd68, 8'd91, 8'd110, 8'd103, 8'd66, 8'd86, 8'd102, 8'd107, 8'd171, 8'd141, 8'd90, 8'd95, 8'd110, 8'd90, 8'd107, 8'd178, 8'd195, 8'd131, 8'd179, 8'd163, 8'd162, 8'd153, 8'd178, 8'd86, 8'd105, 8'd50, 8'd59, 8'd50, 8'd73, 8'd64, 8'd83, 8'd105, 8'd142, 8'd96, 8'd153, 8'd96, 8'd99, 8'd138, 8'd170, 8'd138, 8'd175, 8'd87, 8'd165, 8'd110, 8'd185, 8'd117, 8'd127, 8'd135, 8'd170, 8'd73, 8'd109, 8'd56, 8'd115, 8'd81, 8'd58, 8'd36, 8'd130, 8'd111, 8'd137, 8'd100, 8'd65, 8'd120, 8'd114, 8'd78, 8'd102, 8'd151, 8'd101, 8'd144, 8'd171, 8'd129, 8'd144, 8'd82, 8'd160, 8'd132, 8'd57, 8'd140, 8'd71, 8'd109, 8'd61, 8'd64, 8'd106, 8'd116, 8'd82, 8'd113, 8'd54, 8'd63, 8'd134, 8'd74, 8'd101, 8'd132, 8'd140, 8'd87, 8'd122, 8'd157, 8'd178, 8'd161, 8'd123, 8'd122, 8'd135, 8'd85, 8'd69, 8'd71, 8'd47, 8'd93, 8'd62, 8'd136, 8'd101, 8'd72, 8'd105, 8'd141, 8'd75, 8'd83, 8'd32, 8'd108, 8'd113, 8'd121, 8'd73, 8'd96, 8'd101, 8'd90, 8'd105, 8'd151, 8'd198, 8'd188, 8'd171, 8'd164, 8'd134, 8'd188, 8'd77, 8'd111, 8'd98, 8'd51, 8'd65, 8'd130, 8'd122, 8'd129, 8'd135, 8'd67, 8'd151, 8'd111, 8'd122, 8'd103, 8'd125, 8'd110, 8'd105, 8'd100, 8'd149, 8'd94, 8'd149, 8'd104, 8'd183, 8'd95, 8'd167, 8'd113, 8'd147, 8'd202, 8'd120, 8'd167, 8'd149, 8'd91, 8'd74, 8'd129, 8'd114, 8'd102, 8'd130, 8'd173, 8'd135, 8'd105, 8'd139, 8'd95, 8'd136, 8'd86, 8'd88, 8'd112, 8'd98, 8'd147, 8'd128, 8'd150, 8'd157, 8'd177, 8'd115, 8'd143, 8'd150, 8'd129, 8'd180, 8'd173, 8'd104, 8'd150, 8'd157, 8'd148, 8'd155, 8'd155, 8'd94, 8'd166, 8'd128, 8'd165, 8'd114, 8'd107, 8'd155, 8'd100, 8'd73, 8'd80, 8'd147, 8'd154, 8'd141, 8'd187, 8'd185, 8'd117, 8'd98, 8'd113, 8'd75, 8'd119, 8'd121, 8'd88, 8'd134, 8'd105, 8'd148, 8'd124, 8'd165, 8'd134, 8'd128, 8'd156, 8'd161, 8'd119, 8'd147, 8'd149, 8'd99, 8'd117, 8'd143, 8'd89, 8'd139, 8'd91, 8'd115, 8'd95, 8'd121, 8'd160, 8'd90, 8'd113, 8'd157, 8'd91, 8'd135, 8'd91, 8'd96, 8'd77, 8'd119, 8'd156, 8'd165, 8'd94, 8'd183, 8'd107, 8'd135, 8'd150, 8'd98, 8'd145, 8'd177, 8'd157, 8'd75, 8'd101, 8'd136, 8'd170, 8'd158, 8'd171, 8'd150, 8'd87, 8'd98, 8'd147, 8'd156, 8'd159, 8'd91, 8'd89, 8'd70, 8'd95, 8'd156, 8'd140, 8'd79, 8'd124, 8'd142, 8'd134, 8'd172, 8'd117, 8'd122, 8'd82, 8'd164, 8'd148, 8'd114, 8'd107, 8'd133, 8'd113, 8'd117, 8'd120, 8'd142, 8'd141, 8'd87, 8'd87, 8'd99, 8'd110, 8'd109, 8'd164, 8'd76, 8'd93, 8'd106, 8'd78, 8'd101, 8'd98, 8'd112, 8'd147, 8'd125, 8'd161, 8'd136, 8'd141, 8'd119, 8'd77, 8'd177, 8'd149, 8'd85, 8'd155, 8'd69, 8'd156, 8'd144, 8'd116, 8'd103, 8'd126, 8'd130, 8'd92, 8'd93, 8'd125, 8'd139, 8'd145, 8'd159, 8'd171, 8'd122, 8'd162, 8'd142, 8'd144, 8'd167, 8'd112, 8'd180, 8'd97, 8'd107, 8'd141, 8'd132, 8'd128, 8'd169, 8'd96, 8'd97, 8'd133, 8'd144, 8'd142, 8'd150, 8'd78, 8'd107, 8'd123, 8'd167, 8'd80, 8'd169, 8'd171, 8'd195, 8'd186, 8'd182, 8'd135, 8'd181, 8'd181, 8'd189, 8'd168, 8'd201, 8'd159, 8'd178, 8'd163, 8'd180, 8'd119, 8'd152, 8'd133, 8'd172, 8'd170, 8'd131, 8'd104, 8'd125, 8'd122, 8'd132, 8'd131, 8'd92, 8'd179, 8'd109, 8'd169, 8'd113, 8'd167, 8'd158, 8'd188, 8'd154, 8'd137, 8'd177, 8'd186, 8'd108, 8'd140, 8'd112, 8'd173, 8'd151, 8'd145, 8'd169, 8'd83, 8'd90, 8'd105, 8'd93, 8'd121, 8'd135, 8'd139, 8'd137, 8'd77, 8'd102, 8'd164, 8'd103, 8'd110, 8'd173, 8'd175, 8'd95, 8'd146, 8'd113, 8'd78, 8'd90, 8'd133, 8'd98, 8'd194, 8'd141, 8'd102, 8'd122, 8'd91, 8'd158, 8'd149, 8'd163, 8'd123, 8'd125, 8'd101, 8'd133, 8'd100, 8'd136, 8'd135, 8'd138, 8'd133, 8'd152, 8'd159, 8'd166, 8'd90, 8'd161, 8'd102, 8'd154, 8'd96, 8'd103, 8'd114, 8'd145, 8'd87, 8'd119, 8'd103, 8'd102, 8'd116, 8'd159, 8'd154, 8'd84, 8'd101, 8'd75, 8'd139, 8'd134})
) cell_0_30 (
    .clk(clk),
    .input_index(index_0_29_30),
    .input_value(value_0_29_30),
    .input_result(result_0_29_30),
    .input_enable(enable_0_29_30),
    .output_index(index_0_30_31),
    .output_value(value_0_30_31),
    .output_result(result_0_30_31),
    .output_enable(enable_0_30_31)
);

wire [10-1:0] index_0_31_32;
wire [`DATA_WIDTH-1:0] value_0_31_32;
wire [`DATA_WIDTH*4:0] result_0_31_32;
wire enable_0_31_32;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd156, 8'd105, 8'd94, 8'd153, 8'd133, 8'd132, 8'd69, 8'd156, 8'd153, 8'd138, 8'd55, 8'd59, 8'd72, 8'd65, 8'd55, 8'd78, 8'd87, 8'd93, 8'd95, 8'd153, 8'd121, 8'd131, 8'd145, 8'd146, 8'd83, 8'd112, 8'd124, 8'd98, 8'd99, 8'd115, 8'd112, 8'd90, 8'd73, 8'd120, 8'd153, 8'd176, 8'd136, 8'd105, 8'd146, 8'd92, 8'd143, 8'd115, 8'd172, 8'd127, 8'd85, 8'd82, 8'd186, 8'd117, 8'd89, 8'd98, 8'd112, 8'd92, 8'd171, 8'd79, 8'd136, 8'd73, 8'd103, 8'd158, 8'd139, 8'd93, 8'd179, 8'd166, 8'd188, 8'd145, 8'd94, 8'd99, 8'd89, 8'd137, 8'd138, 8'd141, 8'd124, 8'd101, 8'd125, 8'd139, 8'd125, 8'd109, 8'd129, 8'd96, 8'd102, 8'd160, 8'd98, 8'd116, 8'd167, 8'd118, 8'd108, 8'd75, 8'd61, 8'd127, 8'd155, 8'd112, 8'd117, 8'd95, 8'd145, 8'd167, 8'd142, 8'd88, 8'd135, 8'd78, 8'd121, 8'd81, 8'd69, 8'd99, 8'd128, 8'd111, 8'd105, 8'd106, 8'd139, 8'd101, 8'd119, 8'd128, 8'd94, 8'd124, 8'd102, 8'd135, 8'd154, 8'd155, 8'd81, 8'd95, 8'd116, 8'd178, 8'd157, 8'd105, 8'd94, 8'd96, 8'd95, 8'd120, 8'd70, 8'd148, 8'd80, 8'd131, 8'd161, 8'd91, 8'd149, 8'd110, 8'd164, 8'd81, 8'd152, 8'd157, 8'd86, 8'd127, 8'd101, 8'd104, 8'd113, 8'd153, 8'd93, 8'd114, 8'd85, 8'd103, 8'd138, 8'd146, 8'd77, 8'd162, 8'd89, 8'd70, 8'd115, 8'd101, 8'd121, 8'd89, 8'd164, 8'd172, 8'd127, 8'd80, 8'd141, 8'd159, 8'd116, 8'd115, 8'd89, 8'd165, 8'd148, 8'd149, 8'd68, 8'd149, 8'd89, 8'd130, 8'd133, 8'd87, 8'd71, 8'd116, 8'd120, 8'd112, 8'd141, 8'd97, 8'd125, 8'd79, 8'd127, 8'd57, 8'd134, 8'd137, 8'd156, 8'd165, 8'd94, 8'd135, 8'd149, 8'd85, 8'd105, 8'd111, 8'd95, 8'd79, 8'd95, 8'd61, 8'd113, 8'd63, 8'd90, 8'd156, 8'd57, 8'd138, 8'd97, 8'd87, 8'd85, 8'd78, 8'd84, 8'd34, 8'd102, 8'd46, 8'd58, 8'd112, 8'd112, 8'd130, 8'd101, 8'd109, 8'd108, 8'd104, 8'd62, 8'd140, 8'd100, 8'd151, 8'd60, 8'd76, 8'd104, 8'd48, 8'd96, 8'd91, 8'd115, 8'd56, 8'd146, 8'd147, 8'd66, 8'd60, 8'd87, 8'd77, 8'd98, 8'd98, 8'd74, 8'd68, 8'd116, 8'd101, 8'd158, 8'd94, 8'd156, 8'd102, 8'd90, 8'd76, 8'd104, 8'd136, 8'd82, 8'd29, 8'd84, 8'd49, 8'd145, 8'd61, 8'd77, 8'd85, 8'd114, 8'd90, 8'd165, 8'd73, 8'd65, 8'd109, 8'd69, 8'd126, 8'd134, 8'd112, 8'd81, 8'd92, 8'd153, 8'd85, 8'd90, 8'd100, 8'd92, 8'd98, 8'd129, 8'd118, 8'd13, 8'd102, 8'd81, 8'd126, 8'd74, 8'd155, 8'd67, 8'd149, 8'd67, 8'd84, 8'd134, 8'd151, 8'd63, 8'd98, 8'd96, 8'd111, 8'd112, 8'd72, 8'd143, 8'd130, 8'd87, 8'd142, 8'd126, 8'd97, 8'd150, 8'd108, 8'd71, 8'd115, 8'd57, 8'd117, 8'd87, 8'd69, 8'd84, 8'd71, 8'd79, 8'd103, 8'd137, 8'd152, 8'd124, 8'd95, 8'd61, 8'd65, 8'd98, 8'd48, 8'd57, 8'd99, 8'd137, 8'd105, 8'd94, 8'd76, 8'd151, 8'd64, 8'd159, 8'd163, 8'd89, 8'd65, 8'd102, 8'd71, 8'd47, 8'd133, 8'd58, 8'd80, 8'd149, 8'd77, 8'd175, 8'd165, 8'd102, 8'd142, 8'd128, 8'd103, 8'd64, 8'd59, 8'd145, 8'd125, 8'd138, 8'd129, 8'd164, 8'd122, 8'd170, 8'd73, 8'd80, 8'd95, 8'd92, 8'd68, 8'd63, 8'd63, 8'd49, 8'd58, 8'd128, 8'd83, 8'd115, 8'd156, 8'd109, 8'd147, 8'd147, 8'd160, 8'd104, 8'd110, 8'd63, 8'd73, 8'd149, 8'd102, 8'd126, 8'd114, 8'd130, 8'd127, 8'd172, 8'd105, 8'd105, 8'd117, 8'd101, 8'd144, 8'd83, 8'd85, 8'd104, 8'd116, 8'd156, 8'd96, 8'd113, 8'd124, 8'd99, 8'd126, 8'd164, 8'd193, 8'd136, 8'd68, 8'd111, 8'd159, 8'd103, 8'd134, 8'd145, 8'd147, 8'd115, 8'd101, 8'd88, 8'd102, 8'd120, 8'd143, 8'd89, 8'd139, 8'd77, 8'd62, 8'd108, 8'd91, 8'd130, 8'd166, 8'd96, 8'd98, 8'd93, 8'd144, 8'd213, 8'd177, 8'd121, 8'd132, 8'd115, 8'd91, 8'd134, 8'd150, 8'd96, 8'd133, 8'd151, 8'd157, 8'd83, 8'd94, 8'd64, 8'd159, 8'd101, 8'd159, 8'd108, 8'd85, 8'd80, 8'd50, 8'd112, 8'd139, 8'd105, 8'd95, 8'd86, 8'd183, 8'd184, 8'd167, 8'd84, 8'd119, 8'd154, 8'd90, 8'd155, 8'd119, 8'd178, 8'd91, 8'd130, 8'd70, 8'd60, 8'd84, 8'd89, 8'd149, 8'd152, 8'd125, 8'd193, 8'd145, 8'd95, 8'd116, 8'd150, 8'd87, 8'd133, 8'd83, 8'd171, 8'd159, 8'd113, 8'd112, 8'd75, 8'd117, 8'd116, 8'd73, 8'd103, 8'd100, 8'd125, 8'd145, 8'd61, 8'd142, 8'd105, 8'd125, 8'd146, 8'd97, 8'd86, 8'd124, 8'd115, 8'd153, 8'd131, 8'd123, 8'd99, 8'd119, 8'd164, 8'd165, 8'd128, 8'd97, 8'd186, 8'd124, 8'd123, 8'd164, 8'd110, 8'd77, 8'd123, 8'd158, 8'd66, 8'd112, 8'd72, 8'd100, 8'd98, 8'd118, 8'd95, 8'd86, 8'd142, 8'd151, 8'd171, 8'd158, 8'd155, 8'd79, 8'd133, 8'd155, 8'd125, 8'd181, 8'd122, 8'd151, 8'd158, 8'd176, 8'd147, 8'd112, 8'd88, 8'd121, 8'd66, 8'd120, 8'd98, 8'd113, 8'd95, 8'd80, 8'd49, 8'd55, 8'd68, 8'd123, 8'd105, 8'd137, 8'd177, 8'd168, 8'd138, 8'd127, 8'd146, 8'd148, 8'd183, 8'd147, 8'd171, 8'd100, 8'd112, 8'd92, 8'd167, 8'd126, 8'd112, 8'd124, 8'd55, 8'd52, 8'd53, 8'd99, 8'd87, 8'd99, 8'd67, 8'd50, 8'd143, 8'd93, 8'd127, 8'd125, 8'd163, 8'd156, 8'd110, 8'd136, 8'd156, 8'd77, 8'd92, 8'd78, 8'd96, 8'd129, 8'd126, 8'd76, 8'd171, 8'd153, 8'd141, 8'd99, 8'd73, 8'd92, 8'd88, 8'd127, 8'd146, 8'd56, 8'd138, 8'd139, 8'd116, 8'd142, 8'd147, 8'd154, 8'd74, 8'd76, 8'd77, 8'd119, 8'd76, 8'd125, 8'd106, 8'd95, 8'd100, 8'd80, 8'd117, 8'd137, 8'd154, 8'd142, 8'd76, 8'd101, 8'd89, 8'd104, 8'd74, 8'd60, 8'd134, 8'd133, 8'd80, 8'd164, 8'd86, 8'd163, 8'd157, 8'd146, 8'd111, 8'd146, 8'd155, 8'd122, 8'd122, 8'd65, 8'd50, 8'd109, 8'd116, 8'd46, 8'd52, 8'd103, 8'd56, 8'd104, 8'd65, 8'd122, 8'd55, 8'd100, 8'd48, 8'd61, 8'd157, 8'd129, 8'd167, 8'd80, 8'd133, 8'd102, 8'd121, 8'd127, 8'd160, 8'd77, 8'd132, 8'd135, 8'd53, 8'd123, 8'd50, 8'd38, 8'd98, 8'd46, 8'd97, 8'd71, 8'd99, 8'd77, 8'd91, 8'd14, 8'd106, 8'd69, 8'd76, 8'd103, 8'd127, 8'd124, 8'd151, 8'd122, 8'd75, 8'd91, 8'd158, 8'd162, 8'd67, 8'd149, 8'd62, 8'd46, 8'd130, 8'd110, 8'd105, 8'd37, 8'd65, 8'd117, 8'd84, 8'd39, 8'd69, 8'd74, 8'd37, 8'd34, 8'd73, 8'd122, 8'd55, 8'd54, 8'd137, 8'd103, 8'd76, 8'd115, 8'd95, 8'd110, 8'd136, 8'd114, 8'd79, 8'd94, 8'd104, 8'd119, 8'd94, 8'd60, 8'd90, 8'd92, 8'd114, 8'd116, 8'd97, 8'd78, 8'd131, 8'd83, 8'd82, 8'd134, 8'd94, 8'd72, 8'd147, 8'd106, 8'd148, 8'd95, 8'd103, 8'd142, 8'd72, 8'd78, 8'd98, 8'd72, 8'd130, 8'd92, 8'd88, 8'd125, 8'd82, 8'd139, 8'd158, 8'd107, 8'd142, 8'd114, 8'd83, 8'd137, 8'd145, 8'd147, 8'd141, 8'd114, 8'd152, 8'd81, 8'd159, 8'd82, 8'd81, 8'd143, 8'd146, 8'd97, 8'd142, 8'd71})
) cell_0_31 (
    .clk(clk),
    .input_index(index_0_30_31),
    .input_value(value_0_30_31),
    .input_result(result_0_30_31),
    .input_enable(enable_0_30_31),
    .output_index(index_0_31_32),
    .output_value(value_0_31_32),
    .output_result(result_0_31_32),
    .output_enable(enable_0_31_32)
);

wire [10-1:0] index_0_32_33;
wire [`DATA_WIDTH-1:0] value_0_32_33;
wire [`DATA_WIDTH*4:0] result_0_32_33;
wire enable_0_32_33;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd143, 8'd72, 8'd143, 8'd108, 8'd60, 8'd117, 8'd102, 8'd143, 8'd58, 8'd80, 8'd96, 8'd123, 8'd67, 8'd90, 8'd116, 8'd99, 8'd156, 8'd130, 8'd156, 8'd61, 8'd148, 8'd78, 8'd93, 8'd128, 8'd107, 8'd151, 8'd126, 8'd136, 8'd87, 8'd136, 8'd66, 8'd169, 8'd150, 8'd88, 8'd125, 8'd142, 8'd126, 8'd117, 8'd106, 8'd144, 8'd136, 8'd144, 8'd86, 8'd131, 8'd119, 8'd139, 8'd126, 8'd87, 8'd121, 8'd121, 8'd95, 8'd133, 8'd113, 8'd128, 8'd121, 8'd130, 8'd168, 8'd64, 8'd153, 8'd116, 8'd117, 8'd128, 8'd176, 8'd164, 8'd88, 8'd120, 8'd151, 8'd144, 8'd85, 8'd75, 8'd103, 8'd81, 8'd113, 8'd116, 8'd99, 8'd115, 8'd85, 8'd71, 8'd59, 8'd77, 8'd123, 8'd155, 8'd102, 8'd114, 8'd160, 8'd96, 8'd102, 8'd90, 8'd117, 8'd113, 8'd143, 8'd148, 8'd108, 8'd136, 8'd93, 8'd129, 8'd173, 8'd137, 8'd194, 8'd177, 8'd200, 8'd126, 8'd136, 8'd93, 8'd127, 8'd71, 8'd66, 8'd82, 8'd150, 8'd104, 8'd88, 8'd104, 8'd139, 8'd119, 8'd75, 8'd82, 8'd107, 8'd147, 8'd107, 8'd139, 8'd126, 8'd150, 8'd158, 8'd162, 8'd196, 8'd196, 8'd172, 8'd192, 8'd129, 8'd168, 8'd151, 8'd111, 8'd165, 8'd89, 8'd158, 8'd119, 8'd116, 8'd162, 8'd89, 8'd77, 8'd114, 8'd150, 8'd81, 8'd130, 8'd116, 8'd149, 8'd119, 8'd186, 8'd152, 8'd170, 8'd107, 8'd130, 8'd91, 8'd175, 8'd167, 8'd141, 8'd122, 8'd116, 8'd168, 8'd176, 8'd91, 8'd128, 8'd155, 8'd152, 8'd144, 8'd99, 8'd131, 8'd167, 8'd105, 8'd101, 8'd156, 8'd153, 8'd180, 8'd110, 8'd165, 8'd101, 8'd146, 8'd83, 8'd136, 8'd152, 8'd116, 8'd99, 8'd110, 8'd55, 8'd150, 8'd130, 8'd156, 8'd142, 8'd120, 8'd150, 8'd108, 8'd192, 8'd150, 8'd89, 8'd85, 8'd151, 8'd82, 8'd96, 8'd52, 8'd117, 8'd182, 8'd145, 8'd103, 8'd180, 8'd107, 8'd127, 8'd100, 8'd71, 8'd99, 8'd78, 8'd78, 8'd51, 8'd72, 8'd84, 8'd89, 8'd180, 8'd99, 8'd145, 8'd167, 8'd154, 8'd159, 8'd157, 8'd79, 8'd109, 8'd144, 8'd83, 8'd103, 8'd155, 8'd95, 8'd167, 8'd136, 8'd155, 8'd122, 8'd77, 8'd145, 8'd109, 8'd126, 8'd79, 8'd122, 8'd38, 8'd57, 8'd87, 8'd72, 8'd97, 8'd137, 8'd153, 8'd151, 8'd181, 8'd180, 8'd144, 8'd73, 8'd149, 8'd150, 8'd64, 8'd40, 8'd121, 8'd171, 8'd166, 8'd141, 8'd135, 8'd96, 8'd130, 8'd114, 8'd89, 8'd90, 8'd92, 8'd33, 8'd92, 8'd82, 8'd41, 8'd111, 8'd111, 8'd182, 8'd186, 8'd122, 8'd162, 8'd151, 8'd180, 8'd107, 8'd142, 8'd86, 8'd66, 8'd72, 8'd102, 8'd112, 8'd99, 8'd126, 8'd127, 8'd137, 8'd126, 8'd149, 8'd174, 8'd122, 8'd48, 8'd71, 8'd58, 8'd68, 8'd115, 8'd50, 8'd130, 8'd108, 8'd144, 8'd141, 8'd119, 8'd104, 8'd184, 8'd178, 8'd71, 8'd150, 8'd142, 8'd91, 8'd83, 8'd135, 8'd156, 8'd110, 8'd123, 8'd122, 8'd108, 8'd150, 8'd129, 8'd69, 8'd110, 8'd121, 8'd130, 8'd97, 8'd120, 8'd150, 8'd82, 8'd77, 8'd68, 8'd158, 8'd95, 8'd118, 8'd100, 8'd159, 8'd162, 8'd167, 8'd158, 8'd136, 8'd86, 8'd63, 8'd137, 8'd104, 8'd83, 8'd93, 8'd81, 8'd93, 8'd79, 8'd60, 8'd107, 8'd100, 8'd181, 8'd124, 8'd136, 8'd95, 8'd77, 8'd125, 8'd118, 8'd135, 8'd92, 8'd87, 8'd65, 8'd147, 8'd144, 8'd161, 8'd103, 8'd54, 8'd95, 8'd60, 8'd62, 8'd149, 8'd127, 8'd86, 8'd111, 8'd72, 8'd122, 8'd63, 8'd122, 8'd182, 8'd127, 8'd126, 8'd93, 8'd143, 8'd131, 8'd127, 8'd65, 8'd100, 8'd135, 8'd144, 8'd62, 8'd164, 8'd166, 8'd90, 8'd189, 8'd93, 8'd121, 8'd96, 8'd37, 8'd53, 8'd147, 8'd89, 8'd184, 8'd106, 8'd107, 8'd141, 8'd145, 8'd203, 8'd168, 8'd88, 8'd175, 8'd171, 8'd126, 8'd153, 8'd145, 8'd78, 8'd159, 8'd143, 8'd94, 8'd62, 8'd83, 8'd164, 8'd195, 8'd121, 8'd56, 8'd76, 8'd84, 8'd130, 8'd122, 8'd184, 8'd159, 8'd106, 8'd151, 8'd86, 8'd106, 8'd133, 8'd101, 8'd104, 8'd89, 8'd72, 8'd118, 8'd110, 8'd139, 8'd89, 8'd101, 8'd129, 8'd57, 8'd113, 8'd69, 8'd124, 8'd171, 8'd194, 8'd171, 8'd93, 8'd80, 8'd80, 8'd166, 8'd142, 8'd97, 8'd82, 8'd162, 8'd117, 8'd186, 8'd186, 8'd81, 8'd116, 8'd149, 8'd138, 8'd168, 8'd125, 8'd144, 8'd130, 8'd117, 8'd69, 8'd65, 8'd75, 8'd133, 8'd99, 8'd116, 8'd241, 8'd210, 8'd188, 8'd157, 8'd160, 8'd172, 8'd132, 8'd97, 8'd87, 8'd138, 8'd73, 8'd110, 8'd113, 8'd96, 8'd129, 8'd156, 8'd171, 8'd155, 8'd153, 8'd107, 8'd142, 8'd158, 8'd123, 8'd134, 8'd145, 8'd159, 8'd143, 8'd128, 8'd234, 8'd153, 8'd171, 8'd104, 8'd149, 8'd170, 8'd163, 8'd117, 8'd173, 8'd140, 8'd118, 8'd77, 8'd161, 8'd130, 8'd153, 8'd88, 8'd107, 8'd103, 8'd135, 8'd113, 8'd91, 8'd75, 8'd132, 8'd155, 8'd127, 8'd158, 8'd96, 8'd159, 8'd177, 8'd221, 8'd190, 8'd134, 8'd140, 8'd106, 8'd171, 8'd160, 8'd192, 8'd173, 8'd138, 8'd107, 8'd121, 8'd115, 8'd80, 8'd91, 8'd109, 8'd92, 8'd73, 8'd100, 8'd110, 8'd81, 8'd145, 8'd79, 8'd97, 8'd82, 8'd104, 8'd106, 8'd151, 8'd185, 8'd190, 8'd156, 8'd110, 8'd118, 8'd104, 8'd117, 8'd187, 8'd97, 8'd156, 8'd143, 8'd126, 8'd130, 8'd134, 8'd140, 8'd123, 8'd138, 8'd122, 8'd107, 8'd169, 8'd115, 8'd130, 8'd130, 8'd119, 8'd95, 8'd90, 8'd101, 8'd173, 8'd101, 8'd175, 8'd87, 8'd136, 8'd107, 8'd135, 8'd132, 8'd95, 8'd149, 8'd130, 8'd134, 8'd143, 8'd130, 8'd158, 8'd82, 8'd85, 8'd97, 8'd137, 8'd127, 8'd113, 8'd89, 8'd124, 8'd65, 8'd87, 8'd120, 8'd92, 8'd140, 8'd89, 8'd157, 8'd143, 8'd73, 8'd121, 8'd109, 8'd70, 8'd104, 8'd166, 8'd127, 8'd148, 8'd97, 8'd108, 8'd132, 8'd94, 8'd161, 8'd130, 8'd88, 8'd147, 8'd80, 8'd147, 8'd92, 8'd117, 8'd88, 8'd126, 8'd106, 8'd75, 8'd154, 8'd123, 8'd144, 8'd72, 8'd78, 8'd78, 8'd59, 8'd70, 8'd128, 8'd71, 8'd118, 8'd99, 8'd95, 8'd172, 8'd97, 8'd110, 8'd89, 8'd141, 8'd131, 8'd146, 8'd128, 8'd116, 8'd155, 8'd105, 8'd130, 8'd163, 8'd146, 8'd80, 8'd111, 8'd122, 8'd126, 8'd73, 8'd42, 8'd117, 8'd137, 8'd118, 8'd111, 8'd128, 8'd60, 8'd71, 8'd128, 8'd80, 8'd105, 8'd76, 8'd96, 8'd61, 8'd75, 8'd95, 8'd133, 8'd109, 8'd169, 8'd96, 8'd89, 8'd73, 8'd126, 8'd114, 8'd124, 8'd130, 8'd71, 8'd53, 8'd61, 8'd115, 8'd62, 8'd83, 8'd137, 8'd144, 8'd53, 8'd117, 8'd76, 8'd111, 8'd116, 8'd26, 8'd98, 8'd69, 8'd111, 8'd101, 8'd72, 8'd133, 8'd146, 8'd122, 8'd139, 8'd155, 8'd80, 8'd90, 8'd136, 8'd94, 8'd75, 8'd158, 8'd132, 8'd141, 8'd83, 8'd133, 8'd68, 8'd70, 8'd130, 8'd159, 8'd66, 8'd90, 8'd55, 8'd100, 8'd91, 8'd127, 8'd74, 8'd69, 8'd107, 8'd74, 8'd78, 8'd103, 8'd97, 8'd165, 8'd101, 8'd158, 8'd103, 8'd127, 8'd91, 8'd94, 8'd169, 8'd72, 8'd132, 8'd132, 8'd110, 8'd96, 8'd150, 8'd102, 8'd155, 8'd77, 8'd108, 8'd86, 8'd106, 8'd113, 8'd78, 8'd158, 8'd138, 8'd127, 8'd148, 8'd140, 8'd150, 8'd111, 8'd158})
) cell_0_32 (
    .clk(clk),
    .input_index(index_0_31_32),
    .input_value(value_0_31_32),
    .input_result(result_0_31_32),
    .input_enable(enable_0_31_32),
    .output_index(index_0_32_33),
    .output_value(value_0_32_33),
    .output_result(result_0_32_33),
    .output_enable(enable_0_32_33)
);

wire [10-1:0] index_0_33_34;
wire [`DATA_WIDTH-1:0] value_0_33_34;
wire [`DATA_WIDTH*4:0] result_0_33_34;
wire enable_0_33_34;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd137, 8'd112, 8'd81, 8'd141, 8'd100, 8'd64, 8'd89, 8'd131, 8'd145, 8'd117, 8'd114, 8'd55, 8'd69, 8'd92, 8'd51, 8'd132, 8'd85, 8'd97, 8'd156, 8'd93, 8'd160, 8'd116, 8'd69, 8'd137, 8'd153, 8'd135, 8'd148, 8'd117, 8'd117, 8'd98, 8'd120, 8'd105, 8'd83, 8'd94, 8'd77, 8'd90, 8'd139, 8'd103, 8'd110, 8'd80, 8'd47, 8'd44, 8'd133, 8'd93, 8'd76, 8'd105, 8'd79, 8'd111, 8'd90, 8'd121, 8'd146, 8'd131, 8'd133, 8'd74, 8'd113, 8'd106, 8'd86, 8'd108, 8'd128, 8'd158, 8'd89, 8'd103, 8'd161, 8'd72, 8'd135, 8'd81, 8'd89, 8'd82, 8'd106, 8'd124, 8'd108, 8'd94, 8'd68, 8'd55, 8'd75, 8'd90, 8'd42, 8'd69, 8'd91, 8'd131, 8'd109, 8'd86, 8'd163, 8'd104, 8'd113, 8'd80, 8'd132, 8'd153, 8'd159, 8'd91, 8'd85, 8'd157, 8'd180, 8'd160, 8'd80, 8'd164, 8'd131, 8'd168, 8'd151, 8'd158, 8'd163, 8'd92, 8'd121, 8'd141, 8'd101, 8'd86, 8'd96, 8'd76, 8'd53, 8'd101, 8'd161, 8'd118, 8'd126, 8'd149, 8'd106, 8'd93, 8'd172, 8'd87, 8'd159, 8'd113, 8'd141, 8'd139, 8'd154, 8'd171, 8'd166, 8'd153, 8'd147, 8'd170, 8'd95, 8'd152, 8'd84, 8'd114, 8'd106, 8'd119, 8'd114, 8'd99, 8'd110, 8'd152, 8'd169, 8'd152, 8'd148, 8'd75, 8'd178, 8'd136, 8'd153, 8'd174, 8'd107, 8'd166, 8'd149, 8'd119, 8'd156, 8'd83, 8'd142, 8'd117, 8'd121, 8'd141, 8'd159, 8'd137, 8'd82, 8'd105, 8'd120, 8'd79, 8'd74, 8'd158, 8'd87, 8'd112, 8'd134, 8'd143, 8'd143, 8'd67, 8'd170, 8'd89, 8'd147, 8'd130, 8'd137, 8'd137, 8'd187, 8'd144, 8'd172, 8'd163, 8'd96, 8'd116, 8'd109, 8'd187, 8'd126, 8'd163, 8'd138, 8'd129, 8'd161, 8'd130, 8'd139, 8'd127, 8'd115, 8'd77, 8'd123, 8'd77, 8'd121, 8'd91, 8'd153, 8'd137, 8'd179, 8'd122, 8'd166, 8'd120, 8'd108, 8'd151, 8'd127, 8'd114, 8'd152, 8'd129, 8'd170, 8'd145, 8'd188, 8'd139, 8'd167, 8'd116, 8'd171, 8'd116, 8'd163, 8'd88, 8'd80, 8'd112, 8'd68, 8'd87, 8'd162, 8'd105, 8'd142, 8'd186, 8'd192, 8'd181, 8'd133, 8'd154, 8'd171, 8'd187, 8'd175, 8'd114, 8'd166, 8'd141, 8'd103, 8'd186, 8'd142, 8'd175, 8'd131, 8'd190, 8'd125, 8'd184, 8'd111, 8'd85, 8'd89, 8'd150, 8'd58, 8'd120, 8'd103, 8'd129, 8'd140, 8'd159, 8'd184, 8'd175, 8'd115, 8'd169, 8'd151, 8'd72, 8'd115, 8'd85, 8'd144, 8'd129, 8'd154, 8'd208, 8'd172, 8'd199, 8'd107, 8'd150, 8'd131, 8'd100, 8'd94, 8'd112, 8'd121, 8'd80, 8'd145, 8'd80, 8'd168, 8'd161, 8'd180, 8'd163, 8'd120, 8'd115, 8'd128, 8'd108, 8'd70, 8'd115, 8'd80, 8'd159, 8'd104, 8'd144, 8'd202, 8'd199, 8'd119, 8'd122, 8'd125, 8'd143, 8'd79, 8'd61, 8'd107, 8'd127, 8'd122, 8'd80, 8'd72, 8'd165, 8'd164, 8'd129, 8'd193, 8'd113, 8'd171, 8'd61, 8'd94, 8'd129, 8'd100, 8'd40, 8'd43, 8'd158, 8'd171, 8'd131, 8'd216, 8'd173, 8'd137, 8'd157, 8'd126, 8'd117, 8'd93, 8'd120, 8'd95, 8'd127, 8'd119, 8'd118, 8'd90, 8'd101, 8'd145, 8'd156, 8'd179, 8'd97, 8'd63, 8'd96, 8'd124, 8'd101, 8'd123, 8'd116, 8'd123, 8'd160, 8'd115, 8'd189, 8'd182, 8'd165, 8'd189, 8'd127, 8'd115, 8'd88, 8'd61, 8'd101, 8'd86, 8'd128, 8'd82, 8'd138, 8'd156, 8'd111, 8'd86, 8'd142, 8'd144, 8'd120, 8'd71, 8'd47, 8'd79, 8'd103, 8'd77, 8'd99, 8'd64, 8'd117, 8'd158, 8'd166, 8'd201, 8'd174, 8'd151, 8'd97, 8'd92, 8'd61, 8'd88, 8'd54, 8'd45, 8'd38, 8'd126, 8'd145, 8'd156, 8'd95, 8'd89, 8'd195, 8'd187, 8'd118, 8'd110, 8'd126, 8'd125, 8'd79, 8'd79, 8'd73, 8'd127, 8'd113, 8'd134, 8'd153, 8'd189, 8'd163, 8'd95, 8'd83, 8'd67, 8'd121, 8'd119, 8'd82, 8'd65, 8'd119, 8'd150, 8'd98, 8'd126, 8'd157, 8'd164, 8'd123, 8'd127, 8'd110, 8'd108, 8'd97, 8'd141, 8'd72, 8'd131, 8'd118, 8'd134, 8'd84, 8'd126, 8'd186, 8'd124, 8'd109, 8'd95, 8'd55, 8'd130, 8'd114, 8'd153, 8'd103, 8'd85, 8'd77, 8'd153, 8'd70, 8'd115, 8'd95, 8'd114, 8'd205, 8'd129, 8'd169, 8'd193, 8'd114, 8'd109, 8'd43, 8'd52, 8'd76, 8'd40, 8'd69, 8'd86, 8'd175, 8'd107, 8'd133, 8'd155, 8'd130, 8'd167, 8'd128, 8'd103, 8'd127, 8'd102, 8'd163, 8'd78, 8'd86, 8'd75, 8'd80, 8'd109, 8'd135, 8'd192, 8'd128, 8'd183, 8'd167, 8'd145, 8'd69, 8'd124, 8'd94, 8'd47, 8'd34, 8'd95, 8'd141, 8'd155, 8'd167, 8'd150, 8'd123, 8'd147, 8'd180, 8'd129, 8'd122, 8'd122, 8'd128, 8'd95, 8'd91, 8'd124, 8'd101, 8'd115, 8'd140, 8'd196, 8'd205, 8'd107, 8'd122, 8'd140, 8'd162, 8'd98, 8'd117, 8'd118, 8'd82, 8'd86, 8'd105, 8'd133, 8'd174, 8'd112, 8'd154, 8'd134, 8'd115, 8'd97, 8'd149, 8'd109, 8'd112, 8'd79, 8'd132, 8'd60, 8'd84, 8'd95, 8'd167, 8'd140, 8'd213, 8'd166, 8'd149, 8'd101, 8'd123, 8'd108, 8'd96, 8'd90, 8'd45, 8'd49, 8'd98, 8'd166, 8'd177, 8'd154, 8'd126, 8'd172, 8'd125, 8'd110, 8'd132, 8'd166, 8'd132, 8'd128, 8'd121, 8'd101, 8'd78, 8'd91, 8'd147, 8'd194, 8'd211, 8'd113, 8'd148, 8'd90, 8'd137, 8'd159, 8'd96, 8'd136, 8'd84, 8'd71, 8'd80, 8'd71, 8'd105, 8'd75, 8'd148, 8'd95, 8'd135, 8'd142, 8'd121, 8'd139, 8'd117, 8'd131, 8'd90, 8'd154, 8'd128, 8'd166, 8'd111, 8'd193, 8'd205, 8'd112, 8'd129, 8'd89, 8'd118, 8'd124, 8'd128, 8'd139, 8'd122, 8'd173, 8'd166, 8'd133, 8'd152, 8'd113, 8'd169, 8'd125, 8'd120, 8'd105, 8'd90, 8'd125, 8'd144, 8'd116, 8'd108, 8'd76, 8'd74, 8'd139, 8'd187, 8'd102, 8'd83, 8'd165, 8'd85, 8'd157, 8'd146, 8'd112, 8'd160, 8'd160, 8'd143, 8'd114, 8'd160, 8'd147, 8'd116, 8'd172, 8'd183, 8'd89, 8'd127, 8'd83, 8'd70, 8'd142, 8'd146, 8'd74, 8'd104, 8'd153, 8'd166, 8'd96, 8'd89, 8'd130, 8'd104, 8'd83, 8'd156, 8'd123, 8'd133, 8'd114, 8'd106, 8'd190, 8'd163, 8'd143, 8'd204, 8'd197, 8'd120, 8'd194, 8'd149, 8'd158, 8'd172, 8'd134, 8'd131, 8'd91, 8'd148, 8'd97, 8'd103, 8'd137, 8'd149, 8'd107, 8'd140, 8'd90, 8'd139, 8'd134, 8'd133, 8'd130, 8'd104, 8'd158, 8'd130, 8'd127, 8'd181, 8'd198, 8'd189, 8'd127, 8'd131, 8'd130, 8'd221, 8'd119, 8'd144, 8'd166, 8'd114, 8'd85, 8'd96, 8'd176, 8'd136, 8'd108, 8'd159, 8'd144, 8'd122, 8'd179, 8'd110, 8'd110, 8'd152, 8'd150, 8'd117, 8'd143, 8'd147, 8'd134, 8'd120, 8'd171, 8'd160, 8'd139, 8'd146, 8'd172, 8'd201, 8'd167, 8'd141, 8'd133, 8'd178, 8'd162, 8'd119, 8'd149, 8'd90, 8'd135, 8'd121, 8'd128, 8'd88, 8'd153, 8'd73, 8'd93, 8'd137, 8'd151, 8'd124, 8'd117, 8'd128, 8'd144, 8'd193, 8'd137, 8'd172, 8'd86, 8'd146, 8'd107, 8'd141, 8'd122, 8'd177, 8'd93, 8'd176, 8'd161, 8'd112, 8'd109, 8'd154, 8'd84, 8'd97, 8'd161, 8'd130, 8'd164, 8'd122, 8'd125, 8'd107, 8'd165, 8'd105, 8'd84, 8'd72, 8'd145, 8'd115, 8'd160, 8'd107, 8'd169, 8'd102, 8'd160, 8'd137, 8'd153, 8'd140, 8'd151, 8'd93, 8'd121, 8'd122, 8'd80, 8'd125, 8'd97, 8'd86})
) cell_0_33 (
    .clk(clk),
    .input_index(index_0_32_33),
    .input_value(value_0_32_33),
    .input_result(result_0_32_33),
    .input_enable(enable_0_32_33),
    .output_index(index_0_33_34),
    .output_value(value_0_33_34),
    .output_result(result_0_33_34),
    .output_enable(enable_0_33_34)
);

wire [10-1:0] index_0_34_35;
wire [`DATA_WIDTH-1:0] value_0_34_35;
wire [`DATA_WIDTH*4:0] result_0_34_35;
wire enable_0_34_35;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd75, 8'd128, 8'd134, 8'd102, 8'd176, 8'd105, 8'd169, 8'd160, 8'd129, 8'd174, 8'd147, 8'd150, 8'd165, 8'd102, 8'd154, 8'd145, 8'd158, 8'd131, 8'd177, 8'd173, 8'd92, 8'd149, 8'd125, 8'd124, 8'd150, 8'd156, 8'd100, 8'd148, 8'd108, 8'd83, 8'd125, 8'd82, 8'd82, 8'd132, 8'd123, 8'd165, 8'd165, 8'd202, 8'd174, 8'd186, 8'd172, 8'd148, 8'd212, 8'd145, 8'd169, 8'd207, 8'd151, 8'd216, 8'd144, 8'd111, 8'd128, 8'd127, 8'd122, 8'd74, 8'd115, 8'd128, 8'd152, 8'd146, 8'd149, 8'd135, 8'd157, 8'd100, 8'd173, 8'd188, 8'd147, 8'd131, 8'd181, 8'd144, 8'd156, 8'd106, 8'd152, 8'd116, 8'd194, 8'd154, 8'd148, 8'd124, 8'd169, 8'd170, 8'd133, 8'd122, 8'd117, 8'd114, 8'd162, 8'd129, 8'd132, 8'd67, 8'd75, 8'd128, 8'd126, 8'd172, 8'd100, 8'd93, 8'd141, 8'd166, 8'd138, 8'd152, 8'd116, 8'd99, 8'd136, 8'd111, 8'd148, 8'd116, 8'd86, 8'd83, 8'd91, 8'd102, 8'd99, 8'd78, 8'd121, 8'd154, 8'd80, 8'd110, 8'd118, 8'd159, 8'd119, 8'd76, 8'd125, 8'd169, 8'd134, 8'd105, 8'd157, 8'd168, 8'd143, 8'd82, 8'd126, 8'd164, 8'd68, 8'd89, 8'd139, 8'd111, 8'd124, 8'd147, 8'd163, 8'd154, 8'd95, 8'd120, 8'd134, 8'd154, 8'd164, 8'd94, 8'd122, 8'd159, 8'd145, 8'd150, 8'd155, 8'd141, 8'd85, 8'd91, 8'd117, 8'd117, 8'd83, 8'd148, 8'd156, 8'd116, 8'd106, 8'd115, 8'd82, 8'd77, 8'd131, 8'd162, 8'd122, 8'd121, 8'd175, 8'd145, 8'd138, 8'd126, 8'd139, 8'd121, 8'd82, 8'd119, 8'd88, 8'd159, 8'd58, 8'd79, 8'd103, 8'd102, 8'd70, 8'd148, 8'd129, 8'd154, 8'd70, 8'd150, 8'd111, 8'd84, 8'd100, 8'd90, 8'd76, 8'd158, 8'd120, 8'd124, 8'd136, 8'd141, 8'd114, 8'd104, 8'd103, 8'd152, 8'd84, 8'd62, 8'd155, 8'd108, 8'd129, 8'd153, 8'd116, 8'd140, 8'd107, 8'd140, 8'd135, 8'd79, 8'd106, 8'd158, 8'd135, 8'd140, 8'd142, 8'd57, 8'd142, 8'd80, 8'd129, 8'd117, 8'd83, 8'd62, 8'd97, 8'd119, 8'd82, 8'd100, 8'd133, 8'd115, 8'd132, 8'd116, 8'd111, 8'd138, 8'd93, 8'd138, 8'd116, 8'd132, 8'd123, 8'd73, 8'd152, 8'd137, 8'd128, 8'd87, 8'd147, 8'd93, 8'd65, 8'd154, 8'd128, 8'd91, 8'd129, 8'd67, 8'd128, 8'd119, 8'd114, 8'd161, 8'd86, 8'd103, 8'd83, 8'd106, 8'd134, 8'd87, 8'd79, 8'd102, 8'd99, 8'd87, 8'd64, 8'd98, 8'd128, 8'd124, 8'd122, 8'd126, 8'd128, 8'd100, 8'd81, 8'd134, 8'd132, 8'd151, 8'd84, 8'd95, 8'd114, 8'd168, 8'd92, 8'd92, 8'd105, 8'd120, 8'd77, 8'd108, 8'd138, 8'd98, 8'd72, 8'd145, 8'd103, 8'd93, 8'd68, 8'd110, 8'd149, 8'd97, 8'd188, 8'd148, 8'd86, 8'd118, 8'd111, 8'd55, 8'd52, 8'd93, 8'd111, 8'd67, 8'd85, 8'd75, 8'd142, 8'd91, 8'd103, 8'd97, 8'd63, 8'd136, 8'd82, 8'd67, 8'd122, 8'd150, 8'd145, 8'd86, 8'd82, 8'd96, 8'd92, 8'd113, 8'd124, 8'd135, 8'd77, 8'd97, 8'd87, 8'd125, 8'd107, 8'd64, 8'd141, 8'd102, 8'd173, 8'd98, 8'd112, 8'd161, 8'd89, 8'd101, 8'd104, 8'd129, 8'd82, 8'd134, 8'd148, 8'd67, 8'd150, 8'd83, 8'd119, 8'd173, 8'd111, 8'd119, 8'd148, 8'd92, 8'd61, 8'd109, 8'd84, 8'd138, 8'd58, 8'd86, 8'd134, 8'd77, 8'd150, 8'd130, 8'd93, 8'd108, 8'd60, 8'd49, 8'd127, 8'd87, 8'd113, 8'd90, 8'd76, 8'd125, 8'd156, 8'd109, 8'd179, 8'd128, 8'd196, 8'd130, 8'd112, 8'd126, 8'd61, 8'd117, 8'd126, 8'd110, 8'd131, 8'd66, 8'd103, 8'd158, 8'd149, 8'd148, 8'd120, 8'd123, 8'd94, 8'd79, 8'd97, 8'd110, 8'd119, 8'd69, 8'd91, 8'd137, 8'd127, 8'd121, 8'd102, 8'd173, 8'd194, 8'd171, 8'd151, 8'd80, 8'd98, 8'd116, 8'd112, 8'd124, 8'd155, 8'd136, 8'd92, 8'd176, 8'd172, 8'd164, 8'd134, 8'd140, 8'd138, 8'd156, 8'd58, 8'd51, 8'd91, 8'd91, 8'd158, 8'd151, 8'd151, 8'd86, 8'd162, 8'd106, 8'd143, 8'd169, 8'd108, 8'd62, 8'd95, 8'd155, 8'd104, 8'd144, 8'd121, 8'd106, 8'd190, 8'd164, 8'd104, 8'd142, 8'd103, 8'd151, 8'd160, 8'd73, 8'd129, 8'd53, 8'd91, 8'd103, 8'd69, 8'd138, 8'd77, 8'd131, 8'd113, 8'd183, 8'd178, 8'd214, 8'd152, 8'd104, 8'd165, 8'd153, 8'd129, 8'd171, 8'd163, 8'd179, 8'd135, 8'd185, 8'd121, 8'd134, 8'd114, 8'd140, 8'd139, 8'd70, 8'd73, 8'd124, 8'd83, 8'd124, 8'd104, 8'd154, 8'd115, 8'd69, 8'd83, 8'd177, 8'd130, 8'd147, 8'd175, 8'd106, 8'd173, 8'd125, 8'd134, 8'd139, 8'd113, 8'd110, 8'd140, 8'd103, 8'd146, 8'd107, 8'd162, 8'd121, 8'd89, 8'd108, 8'd129, 8'd70, 8'd128, 8'd142, 8'd94, 8'd128, 8'd110, 8'd95, 8'd145, 8'd149, 8'd184, 8'd156, 8'd148, 8'd108, 8'd153, 8'd105, 8'd177, 8'd130, 8'd94, 8'd149, 8'd138, 8'd95, 8'd109, 8'd155, 8'd131, 8'd130, 8'd131, 8'd98, 8'd132, 8'd62, 8'd118, 8'd104, 8'd77, 8'd141, 8'd116, 8'd160, 8'd162, 8'd120, 8'd147, 8'd149, 8'd130, 8'd166, 8'd130, 8'd141, 8'd94, 8'd134, 8'd170, 8'd78, 8'd157, 8'd129, 8'd146, 8'd142, 8'd161, 8'd71, 8'd129, 8'd149, 8'd121, 8'd97, 8'd129, 8'd97, 8'd142, 8'd139, 8'd148, 8'd102, 8'd103, 8'd183, 8'd140, 8'd119, 8'd162, 8'd97, 8'd117, 8'd98, 8'd146, 8'd93, 8'd164, 8'd93, 8'd116, 8'd161, 8'd100, 8'd100, 8'd119, 8'd128, 8'd141, 8'd118, 8'd86, 8'd68, 8'd111, 8'd57, 8'd137, 8'd97, 8'd134, 8'd91, 8'd143, 8'd141, 8'd102, 8'd95, 8'd142, 8'd151, 8'd154, 8'd131, 8'd131, 8'd67, 8'd144, 8'd86, 8'd152, 8'd119, 8'd160, 8'd95, 8'd80, 8'd93, 8'd105, 8'd80, 8'd102, 8'd106, 8'd156, 8'd93, 8'd88, 8'd88, 8'd100, 8'd77, 8'd49, 8'd113, 8'd96, 8'd103, 8'd150, 8'd77, 8'd141, 8'd118, 8'd141, 8'd66, 8'd103, 8'd85, 8'd130, 8'd60, 8'd140, 8'd110, 8'd151, 8'd71, 8'd150, 8'd134, 8'd154, 8'd147, 8'd137, 8'd79, 8'd103, 8'd130, 8'd166, 8'd114, 8'd137, 8'd114, 8'd91, 8'd109, 8'd119, 8'd103, 8'd72, 8'd95, 8'd88, 8'd117, 8'd78, 8'd78, 8'd124, 8'd153, 8'd106, 8'd94, 8'd109, 8'd137, 8'd80, 8'd128, 8'd144, 8'd124, 8'd155, 8'd151, 8'd130, 8'd84, 8'd126, 8'd158, 8'd86, 8'd80, 8'd104, 8'd146, 8'd149, 8'd122, 8'd125, 8'd145, 8'd147, 8'd121, 8'd81, 8'd114, 8'd161, 8'd109, 8'd164, 8'd152, 8'd165, 8'd150, 8'd119, 8'd166, 8'd100, 8'd86, 8'd116, 8'd152, 8'd83, 8'd156, 8'd97, 8'd139, 8'd136, 8'd113, 8'd97, 8'd115, 8'd143, 8'd130, 8'd98, 8'd104, 8'd93, 8'd107, 8'd178, 8'd144, 8'd75, 8'd124, 8'd149, 8'd85, 8'd87, 8'd120, 8'd162, 8'd161, 8'd110, 8'd118, 8'd161, 8'd107, 8'd110, 8'd114, 8'd110, 8'd125, 8'd64, 8'd89, 8'd73, 8'd153, 8'd84, 8'd138, 8'd129, 8'd106, 8'd152, 8'd163, 8'd145, 8'd168, 8'd131, 8'd160, 8'd154, 8'd82, 8'd122, 8'd120, 8'd74, 8'd160, 8'd154, 8'd97, 8'd152, 8'd170, 8'd113, 8'd153, 8'd142, 8'd113, 8'd166, 8'd116, 8'd69, 8'd76, 8'd128, 8'd149, 8'd161, 8'd144, 8'd106, 8'd125, 8'd108, 8'd135, 8'd128, 8'd150, 8'd134, 8'd144, 8'd123, 8'd76})
) cell_0_34 (
    .clk(clk),
    .input_index(index_0_33_34),
    .input_value(value_0_33_34),
    .input_result(result_0_33_34),
    .input_enable(enable_0_33_34),
    .output_index(index_0_34_35),
    .output_value(value_0_34_35),
    .output_result(result_0_34_35),
    .output_enable(enable_0_34_35)
);

wire [10-1:0] index_0_35_36;
wire [`DATA_WIDTH-1:0] value_0_35_36;
wire [`DATA_WIDTH*4:0] result_0_35_36;
wire enable_0_35_36;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd93, 8'd167, 8'd154, 8'd71, 8'd147, 8'd55, 8'd102, 8'd82, 8'd59, 8'd84, 8'd100, 8'd64, 8'd53, 8'd126, 8'd109, 8'd139, 8'd148, 8'd71, 8'd132, 8'd76, 8'd111, 8'd83, 8'd128, 8'd147, 8'd112, 8'd91, 8'd119, 8'd96, 8'd162, 8'd123, 8'd146, 8'd107, 8'd161, 8'd60, 8'd104, 8'd113, 8'd69, 8'd79, 8'd45, 8'd61, 8'd61, 8'd92, 8'd98, 8'd140, 8'd86, 8'd50, 8'd100, 8'd77, 8'd125, 8'd145, 8'd83, 8'd149, 8'd158, 8'd131, 8'd93, 8'd161, 8'd74, 8'd88, 8'd164, 8'd123, 8'd81, 8'd142, 8'd107, 8'd150, 8'd78, 8'd139, 8'd107, 8'd101, 8'd99, 8'd158, 8'd113, 8'd65, 8'd145, 8'd98, 8'd47, 8'd58, 8'd80, 8'd38, 8'd51, 8'd105, 8'd73, 8'd90, 8'd106, 8'd114, 8'd101, 8'd93, 8'd97, 8'd175, 8'd97, 8'd121, 8'd109, 8'd141, 8'd181, 8'd130, 8'd166, 8'd140, 8'd129, 8'd115, 8'd159, 8'd103, 8'd99, 8'd72, 8'd129, 8'd71, 8'd95, 8'd101, 8'd77, 8'd85, 8'd100, 8'd101, 8'd114, 8'd103, 8'd75, 8'd131, 8'd83, 8'd111, 8'd133, 8'd121, 8'd107, 8'd98, 8'd171, 8'd120, 8'd178, 8'd89, 8'd183, 8'd133, 8'd168, 8'd185, 8'd165, 8'd117, 8'd187, 8'd160, 8'd166, 8'd144, 8'd118, 8'd126, 8'd86, 8'd121, 8'd146, 8'd76, 8'd148, 8'd161, 8'd132, 8'd146, 8'd150, 8'd194, 8'd125, 8'd121, 8'd181, 8'd130, 8'd116, 8'd81, 8'd88, 8'd169, 8'd148, 8'd98, 8'd186, 8'd158, 8'd147, 8'd122, 8'd121, 8'd108, 8'd190, 8'd185, 8'd172, 8'd170, 8'd130, 8'd104, 8'd89, 8'd160, 8'd180, 8'd115, 8'd100, 8'd119, 8'd164, 8'd185, 8'd100, 8'd89, 8'd142, 8'd84, 8'd69, 8'd67, 8'd104, 8'd94, 8'd132, 8'd139, 8'd185, 8'd154, 8'd185, 8'd200, 8'd117, 8'd184, 8'd112, 8'd85, 8'd159, 8'd121, 8'd104, 8'd151, 8'd175, 8'd167, 8'd142, 8'd159, 8'd99, 8'd115, 8'd182, 8'd154, 8'd86, 8'd89, 8'd102, 8'd91, 8'd153, 8'd145, 8'd114, 8'd156, 8'd135, 8'd137, 8'd149, 8'd195, 8'd112, 8'd156, 8'd95, 8'd164, 8'd123, 8'd98, 8'd156, 8'd172, 8'd192, 8'd160, 8'd134, 8'd143, 8'd125, 8'd186, 8'd122, 8'd125, 8'd157, 8'd130, 8'd82, 8'd115, 8'd100, 8'd148, 8'd101, 8'd102, 8'd127, 8'd122, 8'd108, 8'd103, 8'd176, 8'd188, 8'd146, 8'd69, 8'd126, 8'd101, 8'd103, 8'd127, 8'd196, 8'd198, 8'd196, 8'd193, 8'd100, 8'd154, 8'd91, 8'd139, 8'd78, 8'd80, 8'd160, 8'd122, 8'd147, 8'd123, 8'd138, 8'd117, 8'd159, 8'd165, 8'd98, 8'd155, 8'd190, 8'd189, 8'd116, 8'd95, 8'd156, 8'd133, 8'd132, 8'd110, 8'd189, 8'd141, 8'd128, 8'd98, 8'd152, 8'd123, 8'd145, 8'd103, 8'd111, 8'd93, 8'd142, 8'd104, 8'd173, 8'd166, 8'd126, 8'd137, 8'd86, 8'd86, 8'd155, 8'd163, 8'd150, 8'd187, 8'd200, 8'd120, 8'd139, 8'd100, 8'd131, 8'd141, 8'd187, 8'd186, 8'd133, 8'd155, 8'd114, 8'd78, 8'd92, 8'd105, 8'd65, 8'd129, 8'd160, 8'd149, 8'd202, 8'd132, 8'd121, 8'd132, 8'd97, 8'd86, 8'd56, 8'd109, 8'd124, 8'd179, 8'd127, 8'd90, 8'd119, 8'd146, 8'd88, 8'd163, 8'd96, 8'd108, 8'd106, 8'd60, 8'd117, 8'd107, 8'd75, 8'd73, 8'd100, 8'd56, 8'd107, 8'd144, 8'd117, 8'd134, 8'd84, 8'd133, 8'd127, 8'd101, 8'd70, 8'd72, 8'd78, 8'd95, 8'd158, 8'd112, 8'd127, 8'd135, 8'd94, 8'd118, 8'd181, 8'd143, 8'd73, 8'd75, 8'd135, 8'd58, 8'd129, 8'd94, 8'd119, 8'd59, 8'd164, 8'd182, 8'd143, 8'd123, 8'd106, 8'd69, 8'd78, 8'd41, 8'd20, 8'd52, 8'd28, 8'd75, 8'd109, 8'd83, 8'd134, 8'd157, 8'd179, 8'd118, 8'd152, 8'd114, 8'd127, 8'd72, 8'd87, 8'd155, 8'd143, 8'd92, 8'd101, 8'd83, 8'd104, 8'd166, 8'd109, 8'd115, 8'd120, 8'd95, 8'd45, 8'd96, 8'd88, 8'd59, 8'd67, 8'd129, 8'd81, 8'd116, 8'd95, 8'd116, 8'd111, 8'd197, 8'd143, 8'd102, 8'd60, 8'd134, 8'd92, 8'd119, 8'd170, 8'd90, 8'd106, 8'd107, 8'd121, 8'd164, 8'd107, 8'd43, 8'd62, 8'd116, 8'd107, 8'd65, 8'd90, 8'd119, 8'd62, 8'd150, 8'd74, 8'd57, 8'd77, 8'd94, 8'd155, 8'd164, 8'd117, 8'd131, 8'd148, 8'd85, 8'd153, 8'd98, 8'd113, 8'd87, 8'd158, 8'd158, 8'd145, 8'd125, 8'd130, 8'd83, 8'd122, 8'd85, 8'd117, 8'd123, 8'd130, 8'd122, 8'd81, 8'd121, 8'd85, 8'd61, 8'd64, 8'd97, 8'd120, 8'd128, 8'd182, 8'd85, 8'd163, 8'd135, 8'd82, 8'd160, 8'd94, 8'd119, 8'd182, 8'd179, 8'd162, 8'd87, 8'd65, 8'd106, 8'd74, 8'd70, 8'd89, 8'd111, 8'd163, 8'd103, 8'd156, 8'd168, 8'd118, 8'd139, 8'd137, 8'd81, 8'd87, 8'd154, 8'd124, 8'd158, 8'd107, 8'd155, 8'd151, 8'd186, 8'd188, 8'd176, 8'd177, 8'd99, 8'd165, 8'd130, 8'd100, 8'd171, 8'd168, 8'd179, 8'd177, 8'd94, 8'd138, 8'd142, 8'd176, 8'd170, 8'd171, 8'd125, 8'd139, 8'd84, 8'd179, 8'd118, 8'd188, 8'd115, 8'd168, 8'd156, 8'd141, 8'd109, 8'd105, 8'd142, 8'd163, 8'd94, 8'd132, 8'd173, 8'd109, 8'd157, 8'd131, 8'd169, 8'd112, 8'd129, 8'd130, 8'd123, 8'd111, 8'd167, 8'd84, 8'd152, 8'd108, 8'd110, 8'd111, 8'd132, 8'd110, 8'd85, 8'd108, 8'd174, 8'd168, 8'd156, 8'd105, 8'd148, 8'd160, 8'd94, 8'd158, 8'd115, 8'd94, 8'd122, 8'd133, 8'd112, 8'd85, 8'd166, 8'd159, 8'd143, 8'd87, 8'd113, 8'd132, 8'd95, 8'd92, 8'd112, 8'd158, 8'd148, 8'd98, 8'd153, 8'd61, 8'd116, 8'd172, 8'd151, 8'd136, 8'd148, 8'd164, 8'd86, 8'd134, 8'd122, 8'd147, 8'd106, 8'd104, 8'd127, 8'd133, 8'd139, 8'd145, 8'd136, 8'd124, 8'd84, 8'd117, 8'd97, 8'd100, 8'd114, 8'd142, 8'd158, 8'd86, 8'd127, 8'd58, 8'd56, 8'd68, 8'd97, 8'd127, 8'd105, 8'd134, 8'd170, 8'd153, 8'd129, 8'd189, 8'd179, 8'd157, 8'd94, 8'd90, 8'd119, 8'd96, 8'd137, 8'd154, 8'd131, 8'd112, 8'd127, 8'd80, 8'd137, 8'd107, 8'd116, 8'd120, 8'd59, 8'd44, 8'd83, 8'd80, 8'd132, 8'd112, 8'd107, 8'd119, 8'd92, 8'd144, 8'd190, 8'd180, 8'd151, 8'd115, 8'd101, 8'd162, 8'd164, 8'd116, 8'd138, 8'd153, 8'd118, 8'd133, 8'd107, 8'd86, 8'd84, 8'd86, 8'd89, 8'd84, 8'd70, 8'd58, 8'd79, 8'd116, 8'd99, 8'd52, 8'd62, 8'd135, 8'd159, 8'd150, 8'd98, 8'd146, 8'd156, 8'd115, 8'd94, 8'd140, 8'd147, 8'd133, 8'd94, 8'd133, 8'd92, 8'd136, 8'd128, 8'd112, 8'd143, 8'd145, 8'd141, 8'd168, 8'd142, 8'd127, 8'd75, 8'd91, 8'd122, 8'd100, 8'd125, 8'd81, 8'd83, 8'd149, 8'd141, 8'd99, 8'd83, 8'd144, 8'd69, 8'd127, 8'd137, 8'd131, 8'd71, 8'd108, 8'd160, 8'd166, 8'd137, 8'd154, 8'd100, 8'd96, 8'd142, 8'd120, 8'd129, 8'd146, 8'd72, 8'd114, 8'd89, 8'd60, 8'd66, 8'd164, 8'd122, 8'd77, 8'd145, 8'd140, 8'd115, 8'd67, 8'd148, 8'd92, 8'd133, 8'd59, 8'd140, 8'd93, 8'd108, 8'd139, 8'd137, 8'd107, 8'd86, 8'd78, 8'd151, 8'd101, 8'd86, 8'd100, 8'd147, 8'd144, 8'd156, 8'd90, 8'd150, 8'd77, 8'd85, 8'd141, 8'd163, 8'd141, 8'd123, 8'd78, 8'd71, 8'd131, 8'd82, 8'd165, 8'd138, 8'd151, 8'd132, 8'd161, 8'd148, 8'd102, 8'd132})
) cell_0_35 (
    .clk(clk),
    .input_index(index_0_34_35),
    .input_value(value_0_34_35),
    .input_result(result_0_34_35),
    .input_enable(enable_0_34_35),
    .output_index(index_0_35_36),
    .output_value(value_0_35_36),
    .output_result(result_0_35_36),
    .output_enable(enable_0_35_36)
);

wire [10-1:0] index_0_36_37;
wire [`DATA_WIDTH-1:0] value_0_36_37;
wire [`DATA_WIDTH*4:0] result_0_36_37;
wire enable_0_36_37;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd154, 8'd120, 8'd100, 8'd72, 8'd146, 8'd109, 8'd89, 8'd110, 8'd184, 8'd104, 8'd170, 8'd134, 8'd122, 8'd159, 8'd108, 8'd135, 8'd133, 8'd182, 8'd110, 8'd127, 8'd93, 8'd141, 8'd117, 8'd162, 8'd150, 8'd148, 8'd91, 8'd152, 8'd90, 8'd127, 8'd79, 8'd171, 8'd109, 8'd182, 8'd116, 8'd84, 8'd201, 8'd157, 8'd134, 8'd192, 8'd178, 8'd189, 8'd171, 8'd191, 8'd165, 8'd136, 8'd152, 8'd146, 8'd157, 8'd115, 8'd155, 8'd62, 8'd164, 8'd150, 8'd157, 8'd102, 8'd81, 8'd76, 8'd143, 8'd177, 8'd160, 8'd113, 8'd82, 8'd107, 8'd181, 8'd93, 8'd102, 8'd101, 8'd134, 8'd105, 8'd92, 8'd113, 8'd105, 8'd77, 8'd114, 8'd134, 8'd62, 8'd125, 8'd121, 8'd97, 8'd169, 8'd74, 8'd120, 8'd150, 8'd90, 8'd88, 8'd150, 8'd110, 8'd106, 8'd119, 8'd141, 8'd78, 8'd90, 8'd133, 8'd89, 8'd154, 8'd92, 8'd140, 8'd158, 8'd115, 8'd110, 8'd158, 8'd89, 8'd83, 8'd135, 8'd142, 8'd92, 8'd133, 8'd117, 8'd145, 8'd129, 8'd84, 8'd109, 8'd152, 8'd150, 8'd59, 8'd112, 8'd106, 8'd53, 8'd110, 8'd139, 8'd61, 8'd97, 8'd157, 8'd169, 8'd183, 8'd175, 8'd117, 8'd141, 8'd85, 8'd120, 8'd161, 8'd80, 8'd108, 8'd131, 8'd142, 8'd136, 8'd88, 8'd157, 8'd87, 8'd163, 8'd174, 8'd144, 8'd54, 8'd103, 8'd117, 8'd61, 8'd126, 8'd87, 8'd142, 8'd130, 8'd109, 8'd155, 8'd98, 8'd162, 8'd90, 8'd142, 8'd79, 8'd122, 8'd115, 8'd94, 8'd101, 8'd117, 8'd98, 8'd67, 8'd80, 8'd90, 8'd173, 8'd143, 8'd124, 8'd68, 8'd147, 8'd94, 8'd106, 8'd141, 8'd116, 8'd152, 8'd117, 8'd163, 8'd159, 8'd108, 8'd135, 8'd182, 8'd91, 8'd172, 8'd136, 8'd125, 8'd89, 8'd173, 8'd136, 8'd97, 8'd91, 8'd120, 8'd126, 8'd124, 8'd138, 8'd79, 8'd66, 8'd125, 8'd130, 8'd153, 8'd136, 8'd97, 8'd104, 8'd92, 8'd164, 8'd132, 8'd149, 8'd92, 8'd102, 8'd139, 8'd147, 8'd174, 8'd93, 8'd83, 8'd118, 8'd117, 8'd144, 8'd136, 8'd63, 8'd103, 8'd151, 8'd151, 8'd136, 8'd118, 8'd55, 8'd96, 8'd85, 8'd132, 8'd151, 8'd154, 8'd64, 8'd164, 8'd151, 8'd86, 8'd105, 8'd90, 8'd158, 8'd123, 8'd121, 8'd173, 8'd173, 8'd152, 8'd154, 8'd105, 8'd171, 8'd103, 8'd165, 8'd156, 8'd114, 8'd160, 8'd151, 8'd77, 8'd110, 8'd90, 8'd150, 8'd163, 8'd109, 8'd155, 8'd110, 8'd94, 8'd159, 8'd106, 8'd65, 8'd137, 8'd71, 8'd157, 8'd81, 8'd165, 8'd180, 8'd156, 8'd84, 8'd74, 8'd127, 8'd70, 8'd138, 8'd69, 8'd120, 8'd172, 8'd148, 8'd99, 8'd106, 8'd132, 8'd152, 8'd133, 8'd124, 8'd160, 8'd156, 8'd98, 8'd109, 8'd144, 8'd64, 8'd124, 8'd104, 8'd100, 8'd69, 8'd75, 8'd142, 8'd158, 8'd134, 8'd84, 8'd124, 8'd166, 8'd102, 8'd94, 8'd101, 8'd153, 8'd164, 8'd95, 8'd51, 8'd127, 8'd166, 8'd145, 8'd95, 8'd123, 8'd133, 8'd117, 8'd89, 8'd95, 8'd113, 8'd82, 8'd72, 8'd101, 8'd85, 8'd144, 8'd154, 8'd112, 8'd101, 8'd155, 8'd121, 8'd78, 8'd123, 8'd163, 8'd132, 8'd100, 8'd91, 8'd127, 8'd110, 8'd66, 8'd130, 8'd136, 8'd160, 8'd77, 8'd72, 8'd92, 8'd147, 8'd85, 8'd63, 8'd89, 8'd75, 8'd99, 8'd90, 8'd103, 8'd125, 8'd114, 8'd66, 8'd157, 8'd144, 8'd151, 8'd55, 8'd105, 8'd140, 8'd76, 8'd108, 8'd113, 8'd45, 8'd102, 8'd137, 8'd172, 8'd136, 8'd87, 8'd84, 8'd95, 8'd129, 8'd91, 8'd84, 8'd93, 8'd88, 8'd153, 8'd126, 8'd103, 8'd144, 8'd161, 8'd152, 8'd78, 8'd132, 8'd81, 8'd77, 8'd141, 8'd97, 8'd139, 8'd97, 8'd148, 8'd91, 8'd131, 8'd153, 8'd156, 8'd142, 8'd122, 8'd59, 8'd83, 8'd151, 8'd57, 8'd107, 8'd122, 8'd125, 8'd112, 8'd105, 8'd99, 8'd125, 8'd83, 8'd154, 8'd148, 8'd109, 8'd150, 8'd152, 8'd117, 8'd171, 8'd157, 8'd152, 8'd74, 8'd139, 8'd125, 8'd164, 8'd112, 8'd124, 8'd122, 8'd64, 8'd153, 8'd95, 8'd71, 8'd85, 8'd117, 8'd131, 8'd183, 8'd152, 8'd117, 8'd129, 8'd148, 8'd93, 8'd108, 8'd160, 8'd147, 8'd84, 8'd140, 8'd176, 8'd139, 8'd114, 8'd81, 8'd162, 8'd180, 8'd167, 8'd172, 8'd171, 8'd142, 8'd104, 8'd140, 8'd114, 8'd62, 8'd67, 8'd164, 8'd117, 8'd214, 8'd145, 8'd158, 8'd84, 8'd136, 8'd92, 8'd149, 8'd166, 8'd80, 8'd145, 8'd158, 8'd169, 8'd120, 8'd154, 8'd131, 8'd87, 8'd162, 8'd193, 8'd201, 8'd162, 8'd162, 8'd142, 8'd148, 8'd160, 8'd141, 8'd136, 8'd107, 8'd194, 8'd120, 8'd145, 8'd113, 8'd178, 8'd99, 8'd142, 8'd120, 8'd114, 8'd155, 8'd171, 8'd118, 8'd104, 8'd94, 8'd147, 8'd99, 8'd116, 8'd189, 8'd198, 8'd189, 8'd148, 8'd90, 8'd129, 8'd166, 8'd136, 8'd123, 8'd95, 8'd157, 8'd146, 8'd114, 8'd140, 8'd88, 8'd145, 8'd123, 8'd135, 8'd127, 8'd156, 8'd113, 8'd125, 8'd181, 8'd115, 8'd110, 8'd177, 8'd147, 8'd176, 8'd93, 8'd112, 8'd105, 8'd125, 8'd116, 8'd137, 8'd115, 8'd157, 8'd124, 8'd84, 8'd111, 8'd88, 8'd76, 8'd81, 8'd121, 8'd132, 8'd158, 8'd134, 8'd155, 8'd81, 8'd92, 8'd140, 8'd145, 8'd141, 8'd104, 8'd139, 8'd142, 8'd80, 8'd108, 8'd159, 8'd117, 8'd84, 8'd151, 8'd158, 8'd91, 8'd96, 8'd152, 8'd94, 8'd131, 8'd138, 8'd146, 8'd163, 8'd94, 8'd85, 8'd68, 8'd135, 8'd104, 8'd155, 8'd117, 8'd117, 8'd139, 8'd140, 8'd160, 8'd96, 8'd114, 8'd94, 8'd130, 8'd126, 8'd161, 8'd116, 8'd140, 8'd87, 8'd91, 8'd137, 8'd132, 8'd148, 8'd123, 8'd83, 8'd87, 8'd133, 8'd79, 8'd117, 8'd120, 8'd102, 8'd124, 8'd131, 8'd152, 8'd118, 8'd154, 8'd105, 8'd86, 8'd90, 8'd111, 8'd158, 8'd164, 8'd149, 8'd127, 8'd178, 8'd153, 8'd159, 8'd118, 8'd110, 8'd169, 8'd73, 8'd82, 8'd130, 8'd102, 8'd155, 8'd77, 8'd67, 8'd88, 8'd135, 8'd156, 8'd139, 8'd94, 8'd143, 8'd117, 8'd85, 8'd87, 8'd162, 8'd81, 8'd81, 8'd101, 8'd132, 8'd183, 8'd128, 8'd131, 8'd152, 8'd145, 8'd113, 8'd126, 8'd173, 8'd180, 8'd92, 8'd102, 8'd72, 8'd147, 8'd162, 8'd90, 8'd138, 8'd104, 8'd109, 8'd67, 8'd132, 8'd92, 8'd81, 8'd168, 8'd115, 8'd120, 8'd116, 8'd168, 8'd173, 8'd102, 8'd137, 8'd111, 8'd132, 8'd103, 8'd135, 8'd116, 8'd152, 8'd96, 8'd129, 8'd90, 8'd151, 8'd152, 8'd158, 8'd114, 8'd115, 8'd114, 8'd173, 8'd70, 8'd144, 8'd95, 8'd77, 8'd156, 8'd119, 8'd83, 8'd157, 8'd131, 8'd86, 8'd181, 8'd110, 8'd165, 8'd176, 8'd188, 8'd120, 8'd156, 8'd132, 8'd132, 8'd142, 8'd130, 8'd129, 8'd195, 8'd186, 8'd160, 8'd114, 8'd155, 8'd125, 8'd113, 8'd134, 8'd87, 8'd128, 8'd76, 8'd152, 8'd95, 8'd104, 8'd152, 8'd117, 8'd157, 8'd169, 8'd94, 8'd183, 8'd150, 8'd101, 8'd155, 8'd107, 8'd103, 8'd120, 8'd191, 8'd118, 8'd109, 8'd167, 8'd173, 8'd179, 8'd97, 8'd105, 8'd132, 8'd146, 8'd76, 8'd108, 8'd163, 8'd113, 8'd160, 8'd123, 8'd159, 8'd129, 8'd113, 8'd151, 8'd105, 8'd142, 8'd124, 8'd134, 8'd78, 8'd85, 8'd92, 8'd155, 8'd122, 8'd134, 8'd149, 8'd115, 8'd133, 8'd138, 8'd164, 8'd95, 8'd76, 8'd147, 8'd94, 8'd152, 8'd151, 8'd128})
) cell_0_36 (
    .clk(clk),
    .input_index(index_0_35_36),
    .input_value(value_0_35_36),
    .input_result(result_0_35_36),
    .input_enable(enable_0_35_36),
    .output_index(index_0_36_37),
    .output_value(value_0_36_37),
    .output_result(result_0_36_37),
    .output_enable(enable_0_36_37)
);

wire [10-1:0] index_0_37_38;
wire [`DATA_WIDTH-1:0] value_0_37_38;
wire [`DATA_WIDTH*4:0] result_0_37_38;
wire enable_0_37_38;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd161, 8'd117, 8'd162, 8'd77, 8'd77, 8'd83, 8'd115, 8'd154, 8'd152, 8'd102, 8'd152, 8'd94, 8'd86, 8'd160, 8'd75, 8'd154, 8'd95, 8'd158, 8'd110, 8'd118, 8'd119, 8'd103, 8'd160, 8'd70, 8'd150, 8'd75, 8'd139, 8'd112, 8'd110, 8'd153, 8'd123, 8'd113, 8'd89, 8'd161, 8'd98, 8'd138, 8'd138, 8'd182, 8'd178, 8'd138, 8'd155, 8'd120, 8'd186, 8'd183, 8'd176, 8'd148, 8'd189, 8'd148, 8'd184, 8'd105, 8'd91, 8'd162, 8'd157, 8'd152, 8'd157, 8'd166, 8'd129, 8'd145, 8'd136, 8'd98, 8'd102, 8'd131, 8'd128, 8'd148, 8'd153, 8'd144, 8'd182, 8'd149, 8'd149, 8'd111, 8'd166, 8'd167, 8'd121, 8'd97, 8'd120, 8'd89, 8'd84, 8'd91, 8'd108, 8'd150, 8'd133, 8'd93, 8'd169, 8'd101, 8'd117, 8'd148, 8'd121, 8'd125, 8'd141, 8'd186, 8'd158, 8'd94, 8'd96, 8'd110, 8'd149, 8'd150, 8'd154, 8'd148, 8'd145, 8'd159, 8'd103, 8'd137, 8'd124, 8'd81, 8'd97, 8'd55, 8'd143, 8'd48, 8'd49, 8'd140, 8'd139, 8'd144, 8'd154, 8'd152, 8'd141, 8'd170, 8'd189, 8'd129, 8'd138, 8'd116, 8'd78, 8'd104, 8'd58, 8'd140, 8'd158, 8'd107, 8'd112, 8'd91, 8'd100, 8'd105, 8'd125, 8'd75, 8'd116, 8'd64, 8'd69, 8'd50, 8'd108, 8'd76, 8'd132, 8'd124, 8'd163, 8'd140, 8'd98, 8'd140, 8'd95, 8'd150, 8'd151, 8'd113, 8'd127, 8'd131, 8'd142, 8'd110, 8'd156, 8'd91, 8'd97, 8'd173, 8'd73, 8'd68, 8'd88, 8'd172, 8'd94, 8'd96, 8'd155, 8'd70, 8'd91, 8'd119, 8'd163, 8'd163, 8'd115, 8'd125, 8'd101, 8'd134, 8'd155, 8'd112, 8'd156, 8'd73, 8'd85, 8'd136, 8'd85, 8'd118, 8'd104, 8'd80, 8'd117, 8'd87, 8'd90, 8'd111, 8'd150, 8'd152, 8'd149, 8'd75, 8'd84, 8'd79, 8'd99, 8'd136, 8'd94, 8'd85, 8'd116, 8'd95, 8'd119, 8'd126, 8'd123, 8'd88, 8'd92, 8'd113, 8'd81, 8'd69, 8'd150, 8'd131, 8'd123, 8'd81, 8'd124, 8'd100, 8'd162, 8'd109, 8'd142, 8'd76, 8'd78, 8'd143, 8'd92, 8'd99, 8'd118, 8'd135, 8'd152, 8'd107, 8'd102, 8'd84, 8'd166, 8'd146, 8'd135, 8'd106, 8'd64, 8'd63, 8'd80, 8'd114, 8'd141, 8'd60, 8'd82, 8'd78, 8'd166, 8'd146, 8'd101, 8'd107, 8'd162, 8'd135, 8'd115, 8'd67, 8'd141, 8'd50, 8'd78, 8'd63, 8'd98, 8'd140, 8'd127, 8'd179, 8'd145, 8'd157, 8'd156, 8'd147, 8'd72, 8'd131, 8'd144, 8'd145, 8'd132, 8'd153, 8'd120, 8'd83, 8'd170, 8'd195, 8'd190, 8'd186, 8'd168, 8'd115, 8'd153, 8'd91, 8'd54, 8'd78, 8'd55, 8'd110, 8'd93, 8'd129, 8'd130, 8'd188, 8'd128, 8'd113, 8'd102, 8'd88, 8'd112, 8'd78, 8'd149, 8'd101, 8'd153, 8'd94, 8'd112, 8'd166, 8'd175, 8'd162, 8'd133, 8'd123, 8'd153, 8'd154, 8'd76, 8'd155, 8'd104, 8'd147, 8'd86, 8'd103, 8'd113, 8'd124, 8'd176, 8'd125, 8'd117, 8'd140, 8'd84, 8'd94, 8'd64, 8'd79, 8'd107, 8'd151, 8'd83, 8'd151, 8'd163, 8'd111, 8'd105, 8'd167, 8'd120, 8'd165, 8'd97, 8'd120, 8'd144, 8'd128, 8'd144, 8'd90, 8'd153, 8'd72, 8'd153, 8'd115, 8'd158, 8'd143, 8'd194, 8'd160, 8'd114, 8'd141, 8'd128, 8'd100, 8'd117, 8'd91, 8'd174, 8'd75, 8'd92, 8'd88, 8'd99, 8'd121, 8'd71, 8'd100, 8'd152, 8'd163, 8'd69, 8'd92, 8'd122, 8'd160, 8'd147, 8'd123, 8'd90, 8'd113, 8'd93, 8'd194, 8'd126, 8'd71, 8'd118, 8'd157, 8'd155, 8'd164, 8'd86, 8'd70, 8'd88, 8'd148, 8'd138, 8'd131, 8'd143, 8'd147, 8'd127, 8'd105, 8'd88, 8'd147, 8'd135, 8'd99, 8'd93, 8'd109, 8'd88, 8'd125, 8'd110, 8'd71, 8'd118, 8'd122, 8'd177, 8'd167, 8'd149, 8'd178, 8'd165, 8'd182, 8'd123, 8'd105, 8'd151, 8'd110, 8'd111, 8'd49, 8'd59, 8'd91, 8'd89, 8'd93, 8'd96, 8'd148, 8'd122, 8'd130, 8'd152, 8'd170, 8'd162, 8'd142, 8'd147, 8'd120, 8'd117, 8'd140, 8'd84, 8'd131, 8'd139, 8'd159, 8'd185, 8'd124, 8'd125, 8'd149, 8'd116, 8'd130, 8'd99, 8'd144, 8'd88, 8'd84, 8'd140, 8'd138, 8'd151, 8'd85, 8'd149, 8'd96, 8'd96, 8'd167, 8'd71, 8'd76, 8'd78, 8'd166, 8'd135, 8'd132, 8'd118, 8'd121, 8'd126, 8'd112, 8'd94, 8'd173, 8'd142, 8'd100, 8'd98, 8'd149, 8'd119, 8'd87, 8'd97, 8'd158, 8'd83, 8'd151, 8'd107, 8'd136, 8'd101, 8'd131, 8'd167, 8'd160, 8'd88, 8'd134, 8'd106, 8'd137, 8'd139, 8'd85, 8'd66, 8'd141, 8'd119, 8'd151, 8'd140, 8'd77, 8'd127, 8'd83, 8'd130, 8'd90, 8'd54, 8'd134, 8'd73, 8'd106, 8'd124, 8'd130, 8'd185, 8'd151, 8'd104, 8'd106, 8'd151, 8'd156, 8'd94, 8'd93, 8'd158, 8'd86, 8'd101, 8'd112, 8'd144, 8'd110, 8'd130, 8'd99, 8'd108, 8'd147, 8'd98, 8'd83, 8'd98, 8'd81, 8'd85, 8'd120, 8'd162, 8'd135, 8'd153, 8'd181, 8'd128, 8'd123, 8'd108, 8'd72, 8'd74, 8'd130, 8'd152, 8'd157, 8'd160, 8'd95, 8'd75, 8'd92, 8'd157, 8'd166, 8'd118, 8'd133, 8'd82, 8'd137, 8'd92, 8'd128, 8'd113, 8'd83, 8'd120, 8'd153, 8'd91, 8'd169, 8'd124, 8'd109, 8'd172, 8'd135, 8'd152, 8'd130, 8'd121, 8'd77, 8'd76, 8'd152, 8'd108, 8'd127, 8'd92, 8'd118, 8'd68, 8'd163, 8'd147, 8'd86, 8'd166, 8'd151, 8'd104, 8'd96, 8'd156, 8'd157, 8'd91, 8'd138, 8'd153, 8'd146, 8'd171, 8'd145, 8'd129, 8'd98, 8'd163, 8'd87, 8'd72, 8'd61, 8'd105, 8'd79, 8'd63, 8'd72, 8'd137, 8'd117, 8'd157, 8'd145, 8'd97, 8'd143, 8'd89, 8'd155, 8'd152, 8'd98, 8'd134, 8'd156, 8'd139, 8'd134, 8'd106, 8'd176, 8'd122, 8'd129, 8'd119, 8'd109, 8'd124, 8'd92, 8'd64, 8'd103, 8'd117, 8'd163, 8'd141, 8'd71, 8'd164, 8'd83, 8'd117, 8'd114, 8'd133, 8'd113, 8'd142, 8'd77, 8'd162, 8'd124, 8'd153, 8'd81, 8'd78, 8'd71, 8'd138, 8'd90, 8'd132, 8'd143, 8'd87, 8'd73, 8'd152, 8'd135, 8'd64, 8'd125, 8'd113, 8'd149, 8'd142, 8'd152, 8'd121, 8'd155, 8'd173, 8'd104, 8'd137, 8'd145, 8'd110, 8'd169, 8'd164, 8'd153, 8'd131, 8'd158, 8'd76, 8'd106, 8'd130, 8'd132, 8'd82, 8'd87, 8'd132, 8'd145, 8'd110, 8'd65, 8'd74, 8'd54, 8'd118, 8'd117, 8'd130, 8'd119, 8'd127, 8'd126, 8'd157, 8'd131, 8'd173, 8'd184, 8'd101, 8'd91, 8'd168, 8'd111, 8'd158, 8'd92, 8'd78, 8'd130, 8'd129, 8'd74, 8'd93, 8'd153, 8'd140, 8'd132, 8'd100, 8'd117, 8'd123, 8'd142, 8'd118, 8'd140, 8'd120, 8'd134, 8'd119, 8'd72, 8'd174, 8'd148, 8'd88, 8'd136, 8'd129, 8'd114, 8'd124, 8'd153, 8'd96, 8'd142, 8'd108, 8'd116, 8'd110, 8'd88, 8'd180, 8'd101, 8'd193, 8'd94, 8'd185, 8'd110, 8'd97, 8'd158, 8'd153, 8'd129, 8'd141, 8'd146, 8'd141, 8'd133, 8'd83, 8'd169, 8'd118, 8'd74, 8'd148, 8'd156, 8'd95, 8'd101, 8'd140, 8'd140, 8'd97, 8'd122, 8'd104, 8'd93, 8'd131, 8'd149, 8'd175, 8'd166, 8'd172, 8'd129, 8'd81, 8'd106, 8'd152, 8'd148, 8'd71, 8'd75, 8'd99, 8'd109, 8'd131, 8'd142, 8'd143, 8'd168, 8'd77, 8'd127, 8'd155, 8'd136, 8'd151, 8'd132, 8'd169, 8'd146, 8'd169, 8'd175, 8'd129, 8'd92, 8'd158, 8'd116, 8'd162, 8'd117, 8'd132, 8'd93, 8'd96, 8'd89, 8'd106, 8'd148})
) cell_0_37 (
    .clk(clk),
    .input_index(index_0_36_37),
    .input_value(value_0_36_37),
    .input_result(result_0_36_37),
    .input_enable(enable_0_36_37),
    .output_index(index_0_37_38),
    .output_value(value_0_37_38),
    .output_result(result_0_37_38),
    .output_enable(enable_0_37_38)
);

wire [10-1:0] index_0_38_39;
wire [`DATA_WIDTH-1:0] value_0_38_39;
wire [`DATA_WIDTH*4:0] result_0_38_39;
wire enable_0_38_39;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd138, 8'd84, 8'd106, 8'd121, 8'd99, 8'd68, 8'd135, 8'd119, 8'd74, 8'd84, 8'd112, 8'd123, 8'd62, 8'd97, 8'd64, 8'd94, 8'd145, 8'd129, 8'd128, 8'd141, 8'd159, 8'd74, 8'd115, 8'd101, 8'd100, 8'd91, 8'd164, 8'd115, 8'd83, 8'd140, 8'd141, 8'd165, 8'd129, 8'd143, 8'd150, 8'd164, 8'd136, 8'd118, 8'd165, 8'd152, 8'd77, 8'd98, 8'd114, 8'd129, 8'd147, 8'd163, 8'd89, 8'd137, 8'd92, 8'd97, 8'd96, 8'd98, 8'd77, 8'd156, 8'd140, 8'd123, 8'd106, 8'd92, 8'd131, 8'd112, 8'd137, 8'd139, 8'd90, 8'd168, 8'd183, 8'd150, 8'd165, 8'd123, 8'd157, 8'd145, 8'd92, 8'd176, 8'd131, 8'd99, 8'd110, 8'd116, 8'd135, 8'd169, 8'd164, 8'd116, 8'd94, 8'd138, 8'd97, 8'd119, 8'd98, 8'd95, 8'd143, 8'd135, 8'd175, 8'd180, 8'd172, 8'd116, 8'd96, 8'd86, 8'd149, 8'd106, 8'd96, 8'd149, 8'd162, 8'd142, 8'd165, 8'd112, 8'd152, 8'd93, 8'd167, 8'd160, 8'd146, 8'd144, 8'd88, 8'd80, 8'd161, 8'd88, 8'd159, 8'd93, 8'd108, 8'd175, 8'd140, 8'd121, 8'd113, 8'd143, 8'd90, 8'd164, 8'd151, 8'd153, 8'd84, 8'd143, 8'd80, 8'd102, 8'd135, 8'd90, 8'd133, 8'd117, 8'd140, 8'd155, 8'd79, 8'd167, 8'd198, 8'd149, 8'd135, 8'd83, 8'd122, 8'd66, 8'd107, 8'd111, 8'd114, 8'd160, 8'd157, 8'd164, 8'd92, 8'd97, 8'd152, 8'd144, 8'd82, 8'd137, 8'd133, 8'd102, 8'd82, 8'd93, 8'd139, 8'd97, 8'd106, 8'd149, 8'd125, 8'd169, 8'd146, 8'd97, 8'd73, 8'd151, 8'd96, 8'd114, 8'd98, 8'd158, 8'd176, 8'd127, 8'd164, 8'd120, 8'd172, 8'd178, 8'd140, 8'd90, 8'd136, 8'd129, 8'd112, 8'd81, 8'd150, 8'd107, 8'd168, 8'd172, 8'd149, 8'd170, 8'd152, 8'd185, 8'd178, 8'd181, 8'd148, 8'd172, 8'd69, 8'd120, 8'd123, 8'd115, 8'd170, 8'd119, 8'd193, 8'd117, 8'd113, 8'd171, 8'd111, 8'd176, 8'd148, 8'd78, 8'd76, 8'd133, 8'd163, 8'd150, 8'd151, 8'd152, 8'd176, 8'd166, 8'd143, 8'd164, 8'd109, 8'd81, 8'd172, 8'd161, 8'd86, 8'd180, 8'd192, 8'd137, 8'd203, 8'd139, 8'd158, 8'd146, 8'd192, 8'd131, 8'd116, 8'd129, 8'd156, 8'd124, 8'd107, 8'd155, 8'd137, 8'd108, 8'd129, 8'd161, 8'd197, 8'd155, 8'd134, 8'd178, 8'd114, 8'd119, 8'd124, 8'd89, 8'd134, 8'd91, 8'd126, 8'd105, 8'd134, 8'd151, 8'd181, 8'd117, 8'd154, 8'd162, 8'd117, 8'd99, 8'd69, 8'd92, 8'd46, 8'd79, 8'd117, 8'd122, 8'd109, 8'd149, 8'd157, 8'd148, 8'd144, 8'd127, 8'd180, 8'd113, 8'd107, 8'd171, 8'd148, 8'd139, 8'd134, 8'd104, 8'd188, 8'd153, 8'd96, 8'd161, 8'd176, 8'd103, 8'd100, 8'd113, 8'd138, 8'd68, 8'd137, 8'd99, 8'd128, 8'd94, 8'd122, 8'd74, 8'd102, 8'd118, 8'd182, 8'd122, 8'd145, 8'd113, 8'd105, 8'd98, 8'd141, 8'd131, 8'd201, 8'd122, 8'd145, 8'd149, 8'd90, 8'd149, 8'd141, 8'd92, 8'd153, 8'd58, 8'd114, 8'd68, 8'd79, 8'd127, 8'd127, 8'd105, 8'd76, 8'd79, 8'd89, 8'd123, 8'd105, 8'd155, 8'd114, 8'd186, 8'd97, 8'd103, 8'd110, 8'd170, 8'd169, 8'd177, 8'd157, 8'd146, 8'd95, 8'd76, 8'd121, 8'd73, 8'd123, 8'd77, 8'd117, 8'd117, 8'd155, 8'd178, 8'd135, 8'd83, 8'd120, 8'd79, 8'd133, 8'd120, 8'd121, 8'd103, 8'd146, 8'd102, 8'd101, 8'd104, 8'd156, 8'd116, 8'd168, 8'd176, 8'd108, 8'd115, 8'd90, 8'd84, 8'd72, 8'd70, 8'd151, 8'd122, 8'd81, 8'd168, 8'd130, 8'd132, 8'd106, 8'd115, 8'd156, 8'd79, 8'd64, 8'd141, 8'd93, 8'd101, 8'd141, 8'd127, 8'd163, 8'd70, 8'd111, 8'd101, 8'd119, 8'd149, 8'd152, 8'd69, 8'd72, 8'd68, 8'd96, 8'd89, 8'd152, 8'd143, 8'd119, 8'd108, 8'd142, 8'd103, 8'd90, 8'd134, 8'd128, 8'd120, 8'd52, 8'd45, 8'd103, 8'd122, 8'd126, 8'd102, 8'd106, 8'd168, 8'd107, 8'd125, 8'd135, 8'd149, 8'd133, 8'd157, 8'd101, 8'd170, 8'd135, 8'd77, 8'd131, 8'd91, 8'd99, 8'd128, 8'd181, 8'd72, 8'd67, 8'd97, 8'd72, 8'd100, 8'd79, 8'd110, 8'd136, 8'd129, 8'd123, 8'd76, 8'd115, 8'd79, 8'd138, 8'd125, 8'd91, 8'd147, 8'd112, 8'd111, 8'd78, 8'd149, 8'd156, 8'd162, 8'd143, 8'd132, 8'd164, 8'd142, 8'd71, 8'd39, 8'd56, 8'd110, 8'd64, 8'd102, 8'd112, 8'd61, 8'd118, 8'd82, 8'd119, 8'd56, 8'd102, 8'd123, 8'd149, 8'd83, 8'd93, 8'd59, 8'd158, 8'd131, 8'd113, 8'd177, 8'd147, 8'd117, 8'd138, 8'd99, 8'd133, 8'd102, 8'd64, 8'd129, 8'd118, 8'd92, 8'd98, 8'd126, 8'd70, 8'd108, 8'd144, 8'd91, 8'd146, 8'd89, 8'd126, 8'd107, 8'd94, 8'd96, 8'd107, 8'd49, 8'd124, 8'd98, 8'd78, 8'd94, 8'd85, 8'd104, 8'd137, 8'd108, 8'd124, 8'd164, 8'd102, 8'd83, 8'd77, 8'd111, 8'd139, 8'd69, 8'd131, 8'd93, 8'd90, 8'd166, 8'd132, 8'd72, 8'd143, 8'd157, 8'd88, 8'd70, 8'd49, 8'd96, 8'd69, 8'd72, 8'd82, 8'd80, 8'd166, 8'd74, 8'd141, 8'd126, 8'd127, 8'd154, 8'd118, 8'd150, 8'd115, 8'd110, 8'd137, 8'd137, 8'd71, 8'd156, 8'd121, 8'd163, 8'd113, 8'd62, 8'd156, 8'd99, 8'd68, 8'd121, 8'd116, 8'd73, 8'd122, 8'd112, 8'd56, 8'd137, 8'd77, 8'd163, 8'd102, 8'd172, 8'd217, 8'd187, 8'd189, 8'd153, 8'd160, 8'd166, 8'd137, 8'd141, 8'd67, 8'd79, 8'd165, 8'd155, 8'd121, 8'd144, 8'd143, 8'd142, 8'd102, 8'd81, 8'd95, 8'd110, 8'd55, 8'd113, 8'd68, 8'd112, 8'd109, 8'd103, 8'd143, 8'd103, 8'd148, 8'd162, 8'd104, 8'd110, 8'd107, 8'd120, 8'd118, 8'd67, 8'd71, 8'd151, 8'd136, 8'd166, 8'd80, 8'd96, 8'd139, 8'd79, 8'd90, 8'd117, 8'd64, 8'd111, 8'd75, 8'd97, 8'd107, 8'd53, 8'd121, 8'd101, 8'd159, 8'd104, 8'd104, 8'd162, 8'd132, 8'd185, 8'd185, 8'd142, 8'd118, 8'd108, 8'd138, 8'd159, 8'd155, 8'd94, 8'd96, 8'd121, 8'd89, 8'd143, 8'd170, 8'd90, 8'd144, 8'd35, 8'd73, 8'd72, 8'd92, 8'd44, 8'd112, 8'd87, 8'd111, 8'd99, 8'd141, 8'd110, 8'd193, 8'd162, 8'd163, 8'd209, 8'd158, 8'd137, 8'd184, 8'd191, 8'd105, 8'd145, 8'd88, 8'd149, 8'd75, 8'd165, 8'd132, 8'd156, 8'd151, 8'd163, 8'd70, 8'd84, 8'd96, 8'd128, 8'd140, 8'd140, 8'd130, 8'd164, 8'd133, 8'd169, 8'd231, 8'd184, 8'd237, 8'd212, 8'd156, 8'd134, 8'd138, 8'd94, 8'd84, 8'd108, 8'd129, 8'd145, 8'd103, 8'd111, 8'd157, 8'd123, 8'd137, 8'd95, 8'd87, 8'd120, 8'd142, 8'd134, 8'd82, 8'd100, 8'd175, 8'd189, 8'd146, 8'd198, 8'd209, 8'd183, 8'd140, 8'd164, 8'd153, 8'd189, 8'd193, 8'd185, 8'd170, 8'd83, 8'd125, 8'd169, 8'd90, 8'd158, 8'd129, 8'd95, 8'd130, 8'd76, 8'd129, 8'd112, 8'd126, 8'd121, 8'd98, 8'd189, 8'd171, 8'd189, 8'd118, 8'd86, 8'd107, 8'd162, 8'd106, 8'd162, 8'd93, 8'd107, 8'd145, 8'd107, 8'd111, 8'd117, 8'd80, 8'd169, 8'd119, 8'd170, 8'd161, 8'd70, 8'd112, 8'd74, 8'd166, 8'd86, 8'd130, 8'd145, 8'd120, 8'd146, 8'd112, 8'd123, 8'd91, 8'd107, 8'd174, 8'd106, 8'd89, 8'd117, 8'd108, 8'd96, 8'd120, 8'd91, 8'd117, 8'd138, 8'd99, 8'd87, 8'd89, 8'd114})
) cell_0_38 (
    .clk(clk),
    .input_index(index_0_37_38),
    .input_value(value_0_37_38),
    .input_result(result_0_37_38),
    .input_enable(enable_0_37_38),
    .output_index(index_0_38_39),
    .output_value(value_0_38_39),
    .output_result(result_0_38_39),
    .output_enable(enable_0_38_39)
);

wire [10-1:0] index_0_39_40;
wire [`DATA_WIDTH-1:0] value_0_39_40;
wire [`DATA_WIDTH*4:0] result_0_39_40;
wire enable_0_39_40;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd161, 8'd132, 8'd149, 8'd158, 8'd140, 8'd162, 8'd167, 8'd106, 8'd182, 8'd177, 8'd184, 8'd144, 8'd147, 8'd156, 8'd113, 8'd145, 8'd99, 8'd114, 8'd146, 8'd112, 8'd116, 8'd85, 8'd143, 8'd169, 8'd152, 8'd77, 8'd77, 8'd104, 8'd102, 8'd72, 8'd145, 8'd128, 8'd135, 8'd164, 8'd135, 8'd147, 8'd133, 8'd112, 8'd115, 8'd199, 8'd156, 8'd210, 8'd206, 8'd176, 8'd212, 8'd165, 8'd158, 8'd174, 8'd183, 8'd150, 8'd91, 8'd137, 8'd90, 8'd93, 8'd93, 8'd100, 8'd127, 8'd138, 8'd91, 8'd176, 8'd147, 8'd138, 8'd205, 8'd157, 8'd139, 8'd188, 8'd121, 8'd157, 8'd131, 8'd195, 8'd153, 8'd130, 8'd154, 8'd109, 8'd128, 8'd154, 8'd172, 8'd124, 8'd186, 8'd125, 8'd170, 8'd108, 8'd130, 8'd99, 8'd113, 8'd118, 8'd146, 8'd163, 8'd160, 8'd115, 8'd179, 8'd156, 8'd136, 8'd156, 8'd134, 8'd135, 8'd109, 8'd132, 8'd94, 8'd166, 8'd95, 8'd166, 8'd160, 8'd126, 8'd170, 8'd150, 8'd78, 8'd146, 8'd128, 8'd113, 8'd79, 8'd88, 8'd110, 8'd160, 8'd98, 8'd103, 8'd192, 8'd185, 8'd78, 8'd142, 8'd113, 8'd74, 8'd119, 8'd117, 8'd158, 8'd171, 8'd87, 8'd131, 8'd147, 8'd160, 8'd152, 8'd159, 8'd144, 8'd134, 8'd110, 8'd92, 8'd120, 8'd89, 8'd151, 8'd89, 8'd134, 8'd131, 8'd174, 8'd173, 8'd117, 8'd107, 8'd107, 8'd97, 8'd66, 8'd123, 8'd60, 8'd89, 8'd97, 8'd130, 8'd176, 8'd136, 8'd92, 8'd164, 8'd133, 8'd134, 8'd149, 8'd123, 8'd134, 8'd120, 8'd117, 8'd103, 8'd86, 8'd161, 8'd131, 8'd110, 8'd150, 8'd145, 8'd147, 8'd95, 8'd155, 8'd74, 8'd80, 8'd78, 8'd146, 8'd125, 8'd129, 8'd159, 8'd148, 8'd138, 8'd144, 8'd142, 8'd100, 8'd106, 8'd126, 8'd99, 8'd105, 8'd141, 8'd60, 8'd75, 8'd107, 8'd114, 8'd86, 8'd113, 8'd149, 8'd116, 8'd100, 8'd167, 8'd77, 8'd102, 8'd91, 8'd101, 8'd123, 8'd128, 8'd66, 8'd94, 8'd101, 8'd150, 8'd131, 8'd170, 8'd157, 8'd76, 8'd129, 8'd107, 8'd178, 8'd113, 8'd91, 8'd69, 8'd110, 8'd147, 8'd136, 8'd112, 8'd161, 8'd169, 8'd85, 8'd121, 8'd104, 8'd126, 8'd151, 8'd83, 8'd145, 8'd141, 8'd114, 8'd116, 8'd80, 8'd116, 8'd127, 8'd162, 8'd132, 8'd93, 8'd71, 8'd139, 8'd112, 8'd143, 8'd50, 8'd76, 8'd157, 8'd112, 8'd70, 8'd133, 8'd109, 8'd145, 8'd108, 8'd126, 8'd117, 8'd128, 8'd159, 8'd137, 8'd149, 8'd139, 8'd141, 8'd112, 8'd148, 8'd71, 8'd129, 8'd177, 8'd97, 8'd154, 8'd107, 8'd138, 8'd162, 8'd154, 8'd58, 8'd87, 8'd89, 8'd134, 8'd171, 8'd93, 8'd186, 8'd180, 8'd102, 8'd112, 8'd123, 8'd88, 8'd163, 8'd151, 8'd158, 8'd101, 8'd121, 8'd113, 8'd48, 8'd147, 8'd113, 8'd138, 8'd110, 8'd88, 8'd116, 8'd130, 8'd144, 8'd104, 8'd122, 8'd89, 8'd113, 8'd99, 8'd109, 8'd142, 8'd165, 8'd149, 8'd108, 8'd99, 8'd86, 8'd95, 8'd141, 8'd119, 8'd107, 8'd104, 8'd137, 8'd111, 8'd74, 8'd131, 8'd148, 8'd127, 8'd133, 8'd119, 8'd101, 8'd180, 8'd89, 8'd157, 8'd103, 8'd110, 8'd78, 8'd136, 8'd163, 8'd127, 8'd120, 8'd126, 8'd109, 8'd88, 8'd152, 8'd165, 8'd145, 8'd85, 8'd130, 8'd102, 8'd57, 8'd74, 8'd67, 8'd98, 8'd146, 8'd133, 8'd111, 8'd165, 8'd151, 8'd113, 8'd92, 8'd141, 8'd104, 8'd141, 8'd154, 8'd151, 8'd146, 8'd110, 8'd83, 8'd149, 8'd87, 8'd123, 8'd169, 8'd103, 8'd134, 8'd146, 8'd140, 8'd112, 8'd128, 8'd62, 8'd77, 8'd59, 8'd108, 8'd119, 8'd146, 8'd117, 8'd145, 8'd159, 8'd116, 8'd154, 8'd153, 8'd174, 8'd70, 8'd111, 8'd147, 8'd93, 8'd76, 8'd150, 8'd70, 8'd162, 8'd137, 8'd108, 8'd79, 8'd123, 8'd96, 8'd63, 8'd94, 8'd81, 8'd113, 8'd90, 8'd129, 8'd108, 8'd78, 8'd91, 8'd94, 8'd97, 8'd126, 8'd94, 8'd134, 8'd89, 8'd151, 8'd149, 8'd95, 8'd79, 8'd70, 8'd137, 8'd98, 8'd71, 8'd78, 8'd85, 8'd166, 8'd146, 8'd69, 8'd63, 8'd73, 8'd50, 8'd86, 8'd121, 8'd129, 8'd116, 8'd66, 8'd152, 8'd102, 8'd144, 8'd128, 8'd177, 8'd119, 8'd184, 8'd128, 8'd79, 8'd145, 8'd167, 8'd96, 8'd117, 8'd87, 8'd73, 8'd151, 8'd93, 8'd126, 8'd85, 8'd151, 8'd135, 8'd59, 8'd102, 8'd99, 8'd93, 8'd113, 8'd100, 8'd144, 8'd129, 8'd101, 8'd147, 8'd134, 8'd138, 8'd74, 8'd101, 8'd132, 8'd100, 8'd92, 8'd162, 8'd141, 8'd123, 8'd123, 8'd110, 8'd129, 8'd167, 8'd102, 8'd158, 8'd169, 8'd126, 8'd118, 8'd92, 8'd86, 8'd178, 8'd165, 8'd128, 8'd93, 8'd121, 8'd163, 8'd150, 8'd141, 8'd62, 8'd112, 8'd162, 8'd172, 8'd107, 8'd90, 8'd127, 8'd103, 8'd146, 8'd161, 8'd72, 8'd92, 8'd113, 8'd105, 8'd129, 8'd87, 8'd147, 8'd158, 8'd123, 8'd139, 8'd148, 8'd152, 8'd146, 8'd177, 8'd141, 8'd81, 8'd116, 8'd142, 8'd110, 8'd119, 8'd161, 8'd168, 8'd80, 8'd79, 8'd118, 8'd174, 8'd125, 8'd101, 8'd80, 8'd99, 8'd106, 8'd160, 8'd141, 8'd107, 8'd152, 8'd107, 8'd104, 8'd112, 8'd141, 8'd160, 8'd160, 8'd86, 8'd162, 8'd122, 8'd155, 8'd121, 8'd123, 8'd110, 8'd113, 8'd149, 8'd145, 8'd106, 8'd106, 8'd116, 8'd128, 8'd128, 8'd100, 8'd115, 8'd111, 8'd87, 8'd117, 8'd186, 8'd141, 8'd127, 8'd189, 8'd161, 8'd113, 8'd106, 8'd186, 8'd176, 8'd162, 8'd154, 8'd93, 8'd105, 8'd113, 8'd105, 8'd136, 8'd78, 8'd88, 8'd85, 8'd120, 8'd103, 8'd103, 8'd129, 8'd159, 8'd126, 8'd82, 8'd123, 8'd144, 8'd145, 8'd98, 8'd114, 8'd171, 8'd135, 8'd99, 8'd150, 8'd127, 8'd116, 8'd137, 8'd162, 8'd71, 8'd105, 8'd49, 8'd71, 8'd99, 8'd123, 8'd91, 8'd105, 8'd172, 8'd164, 8'd112, 8'd104, 8'd124, 8'd136, 8'd150, 8'd100, 8'd88, 8'd144, 8'd64, 8'd78, 8'd66, 8'd139, 8'd102, 8'd162, 8'd130, 8'd135, 8'd90, 8'd123, 8'd129, 8'd71, 8'd79, 8'd108, 8'd74, 8'd130, 8'd160, 8'd78, 8'd85, 8'd154, 8'd98, 8'd147, 8'd153, 8'd120, 8'd136, 8'd123, 8'd126, 8'd90, 8'd138, 8'd67, 8'd126, 8'd66, 8'd69, 8'd128, 8'd138, 8'd120, 8'd86, 8'd91, 8'd80, 8'd64, 8'd132, 8'd101, 8'd78, 8'd78, 8'd76, 8'd101, 8'd151, 8'd91, 8'd131, 8'd89, 8'd115, 8'd126, 8'd169, 8'd129, 8'd130, 8'd117, 8'd156, 8'd72, 8'd115, 8'd130, 8'd129, 8'd83, 8'd173, 8'd128, 8'd96, 8'd111, 8'd158, 8'd118, 8'd126, 8'd149, 8'd67, 8'd148, 8'd127, 8'd117, 8'd134, 8'd123, 8'd138, 8'd144, 8'd99, 8'd133, 8'd105, 8'd153, 8'd81, 8'd73, 8'd98, 8'd57, 8'd111, 8'd114, 8'd160, 8'd100, 8'd100, 8'd171, 8'd133, 8'd146, 8'd132, 8'd134, 8'd164, 8'd131, 8'd162, 8'd154, 8'd81, 8'd121, 8'd162, 8'd101, 8'd80, 8'd99, 8'd83, 8'd96, 8'd180, 8'd153, 8'd158, 8'd91, 8'd88, 8'd79, 8'd147, 8'd147, 8'd136, 8'd140, 8'd105, 8'd106, 8'd130, 8'd94, 8'd149, 8'd141, 8'd100, 8'd75, 8'd164, 8'd109, 8'd104, 8'd79, 8'd114, 8'd120, 8'd162, 8'd97, 8'd98, 8'd151, 8'd145, 8'd96, 8'd99, 8'd105, 8'd155, 8'd73, 8'd172, 8'd103, 8'd131, 8'd88, 8'd99, 8'd146, 8'd124, 8'd98, 8'd107, 8'd110, 8'd109, 8'd107, 8'd123, 8'd144, 8'd95})
) cell_0_39 (
    .clk(clk),
    .input_index(index_0_38_39),
    .input_value(value_0_38_39),
    .input_result(result_0_38_39),
    .input_enable(enable_0_38_39),
    .output_index(index_0_39_40),
    .output_value(value_0_39_40),
    .output_result(result_0_39_40),
    .output_enable(enable_0_39_40)
);

wire [10-1:0] index_0_40_41;
wire [`DATA_WIDTH-1:0] value_0_40_41;
wire [`DATA_WIDTH*4:0] result_0_40_41;
wire enable_0_40_41;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd102, 8'd144, 8'd141, 8'd127, 8'd156, 8'd126, 8'd119, 8'd99, 8'd93, 8'd116, 8'd110, 8'd119, 8'd143, 8'd164, 8'd157, 8'd172, 8'd123, 8'd108, 8'd103, 8'd116, 8'd98, 8'd86, 8'd137, 8'd80, 8'd78, 8'd94, 8'd86, 8'd150, 8'd74, 8'd144, 8'd149, 8'd86, 8'd109, 8'd91, 8'd124, 8'd87, 8'd169, 8'd194, 8'd169, 8'd195, 8'd150, 8'd193, 8'd160, 8'd131, 8'd110, 8'd184, 8'd187, 8'd123, 8'd132, 8'd116, 8'd94, 8'd141, 8'd87, 8'd151, 8'd86, 8'd132, 8'd131, 8'd131, 8'd111, 8'd71, 8'd104, 8'd103, 8'd102, 8'd184, 8'd96, 8'd129, 8'd115, 8'd83, 8'd100, 8'd87, 8'd90, 8'd102, 8'd106, 8'd82, 8'd130, 8'd136, 8'd122, 8'd123, 8'd137, 8'd154, 8'd90, 8'd97, 8'd121, 8'd71, 8'd71, 8'd117, 8'd61, 8'd74, 8'd92, 8'd104, 8'd70, 8'd75, 8'd128, 8'd95, 8'd114, 8'd116, 8'd96, 8'd99, 8'd93, 8'd114, 8'd114, 8'd170, 8'd178, 8'd150, 8'd141, 8'd153, 8'd105, 8'd145, 8'd163, 8'd89, 8'd148, 8'd123, 8'd101, 8'd166, 8'd127, 8'd74, 8'd57, 8'd131, 8'd152, 8'd74, 8'd133, 8'd80, 8'd181, 8'd187, 8'd154, 8'd114, 8'd120, 8'd119, 8'd152, 8'd173, 8'd133, 8'd173, 8'd93, 8'd129, 8'd114, 8'd112, 8'd148, 8'd99, 8'd89, 8'd140, 8'd99, 8'd103, 8'd97, 8'd60, 8'd62, 8'd74, 8'd115, 8'd125, 8'd135, 8'd75, 8'd133, 8'd95, 8'd121, 8'd183, 8'd78, 8'd140, 8'd99, 8'd168, 8'd74, 8'd157, 8'd166, 8'd126, 8'd132, 8'd69, 8'd84, 8'd113, 8'd109, 8'd147, 8'd79, 8'd77, 8'd55, 8'd58, 8'd59, 8'd61, 8'd81, 8'd133, 8'd116, 8'd146, 8'd112, 8'd95, 8'd100, 8'd103, 8'd125, 8'd144, 8'd142, 8'd129, 8'd104, 8'd157, 8'd174, 8'd95, 8'd87, 8'd130, 8'd65, 8'd103, 8'd147, 8'd101, 8'd89, 8'd76, 8'd60, 8'd136, 8'd75, 8'd135, 8'd117, 8'd108, 8'd118, 8'd68, 8'd109, 8'd123, 8'd81, 8'd65, 8'd123, 8'd71, 8'd71, 8'd75, 8'd111, 8'd119, 8'd102, 8'd80, 8'd138, 8'd111, 8'd74, 8'd125, 8'd166, 8'd79, 8'd100, 8'd100, 8'd118, 8'd79, 8'd70, 8'd62, 8'd140, 8'd117, 8'd114, 8'd160, 8'd78, 8'd87, 8'd144, 8'd93, 8'd59, 8'd129, 8'd61, 8'd79, 8'd91, 8'd138, 8'd89, 8'd72, 8'd104, 8'd110, 8'd94, 8'd81, 8'd161, 8'd173, 8'd141, 8'd101, 8'd83, 8'd92, 8'd108, 8'd79, 8'd116, 8'd128, 8'd82, 8'd148, 8'd69, 8'd144, 8'd83, 8'd62, 8'd111, 8'd95, 8'd79, 8'd120, 8'd69, 8'd162, 8'd71, 8'd74, 8'd116, 8'd107, 8'd111, 8'd96, 8'd118, 8'd161, 8'd118, 8'd90, 8'd29, 8'd129, 8'd137, 8'd112, 8'd138, 8'd139, 8'd139, 8'd64, 8'd118, 8'd126, 8'd139, 8'd95, 8'd96, 8'd128, 8'd92, 8'd141, 8'd109, 8'd128, 8'd73, 8'd112, 8'd96, 8'd162, 8'd71, 8'd92, 8'd159, 8'd119, 8'd116, 8'd113, 8'd104, 8'd110, 8'd106, 8'd124, 8'd157, 8'd93, 8'd145, 8'd64, 8'd114, 8'd107, 8'd87, 8'd78, 8'd96, 8'd79, 8'd106, 8'd94, 8'd162, 8'd95, 8'd164, 8'd112, 8'd144, 8'd168, 8'd123, 8'd125, 8'd173, 8'd155, 8'd64, 8'd103, 8'd93, 8'd136, 8'd153, 8'd161, 8'd119, 8'd140, 8'd152, 8'd126, 8'd163, 8'd121, 8'd67, 8'd137, 8'd156, 8'd81, 8'd133, 8'd105, 8'd145, 8'd100, 8'd138, 8'd105, 8'd80, 8'd103, 8'd102, 8'd99, 8'd87, 8'd85, 8'd149, 8'd60, 8'd49, 8'd109, 8'd130, 8'd82, 8'd154, 8'd68, 8'd147, 8'd88, 8'd92, 8'd82, 8'd172, 8'd108, 8'd127, 8'd138, 8'd63, 8'd149, 8'd162, 8'd94, 8'd122, 8'd107, 8'd141, 8'd173, 8'd90, 8'd161, 8'd141, 8'd107, 8'd143, 8'd67, 8'd60, 8'd147, 8'd121, 8'd150, 8'd156, 8'd103, 8'd140, 8'd115, 8'd148, 8'd158, 8'd170, 8'd173, 8'd142, 8'd150, 8'd119, 8'd75, 8'd119, 8'd123, 8'd171, 8'd124, 8'd148, 8'd134, 8'd104, 8'd111, 8'd180, 8'd132, 8'd150, 8'd55, 8'd91, 8'd167, 8'd171, 8'd103, 8'd181, 8'd92, 8'd126, 8'd139, 8'd185, 8'd172, 8'd121, 8'd143, 8'd196, 8'd147, 8'd149, 8'd178, 8'd142, 8'd106, 8'd119, 8'd175, 8'd143, 8'd160, 8'd176, 8'd94, 8'd116, 8'd157, 8'd125, 8'd101, 8'd128, 8'd135, 8'd119, 8'd121, 8'd117, 8'd112, 8'd102, 8'd107, 8'd142, 8'd173, 8'd95, 8'd147, 8'd138, 8'd153, 8'd111, 8'd163, 8'd156, 8'd187, 8'd155, 8'd105, 8'd172, 8'd131, 8'd87, 8'd166, 8'd148, 8'd84, 8'd174, 8'd87, 8'd65, 8'd133, 8'd108, 8'd126, 8'd90, 8'd131, 8'd120, 8'd127, 8'd118, 8'd180, 8'd159, 8'd153, 8'd117, 8'd117, 8'd127, 8'd159, 8'd146, 8'd122, 8'd160, 8'd174, 8'd115, 8'd122, 8'd87, 8'd94, 8'd168, 8'd96, 8'd104, 8'd106, 8'd72, 8'd125, 8'd94, 8'd109, 8'd91, 8'd175, 8'd153, 8'd145, 8'd91, 8'd126, 8'd153, 8'd125, 8'd70, 8'd107, 8'd113, 8'd124, 8'd153, 8'd80, 8'd123, 8'd103, 8'd110, 8'd127, 8'd127, 8'd101, 8'd85, 8'd113, 8'd152, 8'd79, 8'd137, 8'd128, 8'd120, 8'd127, 8'd107, 8'd99, 8'd102, 8'd122, 8'd119, 8'd110, 8'd102, 8'd121, 8'd142, 8'd101, 8'd59, 8'd139, 8'd150, 8'd70, 8'd84, 8'd81, 8'd90, 8'd122, 8'd119, 8'd125, 8'd94, 8'd133, 8'd145, 8'd144, 8'd62, 8'd102, 8'd104, 8'd149, 8'd88, 8'd160, 8'd167, 8'd179, 8'd144, 8'd145, 8'd156, 8'd129, 8'd161, 8'd157, 8'd102, 8'd130, 8'd79, 8'd65, 8'd161, 8'd166, 8'd128, 8'd129, 8'd91, 8'd135, 8'd74, 8'd126, 8'd77, 8'd99, 8'd154, 8'd109, 8'd128, 8'd153, 8'd148, 8'd131, 8'd143, 8'd158, 8'd157, 8'd116, 8'd154, 8'd161, 8'd161, 8'd72, 8'd115, 8'd157, 8'd154, 8'd137, 8'd152, 8'd140, 8'd93, 8'd70, 8'd174, 8'd164, 8'd83, 8'd76, 8'd139, 8'd154, 8'd120, 8'd147, 8'd68, 8'd90, 8'd92, 8'd132, 8'd68, 8'd144, 8'd108, 8'd91, 8'd66, 8'd161, 8'd98, 8'd71, 8'd149, 8'd156, 8'd109, 8'd138, 8'd160, 8'd118, 8'd129, 8'd164, 8'd97, 8'd81, 8'd152, 8'd91, 8'd118, 8'd148, 8'd86, 8'd72, 8'd156, 8'd95, 8'd134, 8'd158, 8'd139, 8'd115, 8'd108, 8'd61, 8'd113, 8'd142, 8'd158, 8'd103, 8'd94, 8'd113, 8'd153, 8'd93, 8'd71, 8'd162, 8'd128, 8'd95, 8'd88, 8'd137, 8'd169, 8'd103, 8'd127, 8'd122, 8'd132, 8'd155, 8'd137, 8'd74, 8'd124, 8'd60, 8'd74, 8'd100, 8'd76, 8'd121, 8'd94, 8'd135, 8'd141, 8'd142, 8'd65, 8'd113, 8'd56, 8'd124, 8'd164, 8'd83, 8'd138, 8'd145, 8'd124, 8'd174, 8'd118, 8'd151, 8'd141, 8'd147, 8'd124, 8'd163, 8'd175, 8'd84, 8'd135, 8'd140, 8'd114, 8'd113, 8'd73, 8'd114, 8'd102, 8'd72, 8'd128, 8'd167, 8'd94, 8'd168, 8'd109, 8'd161, 8'd104, 8'd113, 8'd162, 8'd163, 8'd147, 8'd85, 8'd160, 8'd149, 8'd80, 8'd91, 8'd129, 8'd162, 8'd157, 8'd138, 8'd163, 8'd174, 8'd102, 8'd125, 8'd138, 8'd69, 8'd125, 8'd106, 8'd119, 8'd133, 8'd128, 8'd90, 8'd89, 8'd108, 8'd147, 8'd98, 8'd104, 8'd148, 8'd169, 8'd148, 8'd96, 8'd100, 8'd132, 8'd142, 8'd81, 8'd106, 8'd87, 8'd117, 8'd110, 8'd87, 8'd120, 8'd170, 8'd77, 8'd161, 8'd74, 8'd102, 8'd172, 8'd74, 8'd154, 8'd113, 8'd117, 8'd123, 8'd109, 8'd161, 8'd149, 8'd160, 8'd121, 8'd142, 8'd113, 8'd143})
) cell_0_40 (
    .clk(clk),
    .input_index(index_0_39_40),
    .input_value(value_0_39_40),
    .input_result(result_0_39_40),
    .input_enable(enable_0_39_40),
    .output_index(index_0_40_41),
    .output_value(value_0_40_41),
    .output_result(result_0_40_41),
    .output_enable(enable_0_40_41)
);

wire [10-1:0] index_0_41_42;
wire [`DATA_WIDTH-1:0] value_0_41_42;
wire [`DATA_WIDTH*4:0] result_0_41_42;
wire enable_0_41_42;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd109, 8'd85, 8'd127, 8'd159, 8'd129, 8'd86, 8'd103, 8'd98, 8'd158, 8'd148, 8'd109, 8'd105, 8'd113, 8'd196, 8'd146, 8'd109, 8'd93, 8'd108, 8'd100, 8'd124, 8'd155, 8'd109, 8'd133, 8'd146, 8'd118, 8'd146, 8'd111, 8'd122, 8'd132, 8'd78, 8'd147, 8'd150, 8'd164, 8'd133, 8'd149, 8'd119, 8'd160, 8'd197, 8'd161, 8'd171, 8'd171, 8'd129, 8'd183, 8'd115, 8'd128, 8'd109, 8'd119, 8'd118, 8'd129, 8'd110, 8'd131, 8'd121, 8'd153, 8'd75, 8'd131, 8'd105, 8'd166, 8'd155, 8'd114, 8'd90, 8'd115, 8'd122, 8'd163, 8'd116, 8'd99, 8'd181, 8'd134, 8'd169, 8'd150, 8'd145, 8'd172, 8'd113, 8'd160, 8'd186, 8'd131, 8'd196, 8'd187, 8'd154, 8'd132, 8'd109, 8'd82, 8'd122, 8'd114, 8'd120, 8'd145, 8'd165, 8'd82, 8'd114, 8'd100, 8'd115, 8'd159, 8'd134, 8'd90, 8'd79, 8'd95, 8'd154, 8'd142, 8'd158, 8'd157, 8'd125, 8'd135, 8'd164, 8'd130, 8'd174, 8'd128, 8'd175, 8'd152, 8'd152, 8'd160, 8'd126, 8'd168, 8'd157, 8'd147, 8'd112, 8'd58, 8'd148, 8'd120, 8'd118, 8'd121, 8'd142, 8'd60, 8'd118, 8'd138, 8'd102, 8'd107, 8'd126, 8'd110, 8'd98, 8'd105, 8'd138, 8'd162, 8'd164, 8'd147, 8'd133, 8'd139, 8'd119, 8'd90, 8'd153, 8'd151, 8'd93, 8'd101, 8'd154, 8'd132, 8'd86, 8'd87, 8'd66, 8'd148, 8'd85, 8'd138, 8'd71, 8'd83, 8'd107, 8'd96, 8'd82, 8'd96, 8'd92, 8'd113, 8'd163, 8'd86, 8'd110, 8'd87, 8'd94, 8'd125, 8'd58, 8'd141, 8'd102, 8'd149, 8'd82, 8'd149, 8'd126, 8'd120, 8'd110, 8'd91, 8'd54, 8'd74, 8'd114, 8'd81, 8'd113, 8'd130, 8'd80, 8'd140, 8'd154, 8'd82, 8'd70, 8'd126, 8'd88, 8'd157, 8'd93, 8'd165, 8'd123, 8'd87, 8'd139, 8'd134, 8'd80, 8'd110, 8'd163, 8'd146, 8'd101, 8'd123, 8'd90, 8'd119, 8'd119, 8'd93, 8'd130, 8'd123, 8'd98, 8'd58, 8'd80, 8'd90, 8'd118, 8'd103, 8'd134, 8'd115, 8'd118, 8'd67, 8'd105, 8'd105, 8'd138, 8'd131, 8'd126, 8'd134, 8'd79, 8'd162, 8'd152, 8'd159, 8'd101, 8'd135, 8'd89, 8'd79, 8'd52, 8'd90, 8'd133, 8'd97, 8'd79, 8'd123, 8'd114, 8'd124, 8'd64, 8'd86, 8'd135, 8'd74, 8'd115, 8'd72, 8'd110, 8'd145, 8'd102, 8'd95, 8'd146, 8'd108, 8'd81, 8'd169, 8'd149, 8'd83, 8'd111, 8'd57, 8'd51, 8'd63, 8'd113, 8'd51, 8'd135, 8'd88, 8'd80, 8'd63, 8'd54, 8'd147, 8'd121, 8'd73, 8'd130, 8'd92, 8'd145, 8'd65, 8'd118, 8'd139, 8'd56, 8'd149, 8'd161, 8'd130, 8'd120, 8'd150, 8'd140, 8'd108, 8'd153, 8'd75, 8'd95, 8'd66, 8'd80, 8'd111, 8'd154, 8'd81, 8'd136, 8'd148, 8'd145, 8'd139, 8'd104, 8'd66, 8'd83, 8'd115, 8'd90, 8'd153, 8'd106, 8'd140, 8'd126, 8'd109, 8'd108, 8'd73, 8'd171, 8'd92, 8'd97, 8'd133, 8'd120, 8'd28, 8'd77, 8'd62, 8'd76, 8'd129, 8'd146, 8'd143, 8'd169, 8'd136, 8'd152, 8'd135, 8'd70, 8'd134, 8'd58, 8'd72, 8'd88, 8'd65, 8'd109, 8'd139, 8'd129, 8'd85, 8'd157, 8'd163, 8'd125, 8'd129, 8'd99, 8'd79, 8'd59, 8'd139, 8'd123, 8'd132, 8'd101, 8'd128, 8'd93, 8'd87, 8'd156, 8'd138, 8'd136, 8'd160, 8'd83, 8'd109, 8'd110, 8'd51, 8'd108, 8'd116, 8'd76, 8'd117, 8'd93, 8'd110, 8'd106, 8'd101, 8'd123, 8'd88, 8'd160, 8'd144, 8'd130, 8'd129, 8'd148, 8'd132, 8'd139, 8'd117, 8'd149, 8'd136, 8'd103, 8'd130, 8'd115, 8'd124, 8'd140, 8'd55, 8'd99, 8'd49, 8'd88, 8'd61, 8'd127, 8'd124, 8'd160, 8'd182, 8'd178, 8'd177, 8'd119, 8'd141, 8'd136, 8'd97, 8'd51, 8'd111, 8'd101, 8'd155, 8'd134, 8'd76, 8'd90, 8'd158, 8'd117, 8'd159, 8'd105, 8'd145, 8'd89, 8'd67, 8'd93, 8'd58, 8'd123, 8'd78, 8'd129, 8'd95, 8'd91, 8'd171, 8'd159, 8'd200, 8'd191, 8'd158, 8'd131, 8'd110, 8'd139, 8'd93, 8'd115, 8'd124, 8'd174, 8'd136, 8'd167, 8'd187, 8'd105, 8'd128, 8'd108, 8'd118, 8'd94, 8'd132, 8'd104, 8'd68, 8'd83, 8'd128, 8'd178, 8'd175, 8'd100, 8'd184, 8'd114, 8'd116, 8'd130, 8'd184, 8'd105, 8'd79, 8'd79, 8'd96, 8'd127, 8'd150, 8'd105, 8'd154, 8'd177, 8'd104, 8'd117, 8'd116, 8'd133, 8'd152, 8'd160, 8'd153, 8'd101, 8'd82, 8'd78, 8'd101, 8'd85, 8'd94, 8'd149, 8'd183, 8'd94, 8'd151, 8'd108, 8'd130, 8'd110, 8'd163, 8'd43, 8'd63, 8'd80, 8'd148, 8'd144, 8'd128, 8'd105, 8'd155, 8'd127, 8'd191, 8'd166, 8'd187, 8'd110, 8'd109, 8'd120, 8'd167, 8'd77, 8'd76, 8'd166, 8'd127, 8'd157, 8'd90, 8'd120, 8'd168, 8'd142, 8'd145, 8'd94, 8'd90, 8'd82, 8'd103, 8'd60, 8'd128, 8'd158, 8'd129, 8'd90, 8'd146, 8'd170, 8'd137, 8'd197, 8'd154, 8'd98, 8'd97, 8'd81, 8'd160, 8'd124, 8'd148, 8'd106, 8'd108, 8'd138, 8'd107, 8'd132, 8'd144, 8'd155, 8'd138, 8'd143, 8'd121, 8'd61, 8'd115, 8'd132, 8'd107, 8'd113, 8'd153, 8'd180, 8'd122, 8'd151, 8'd164, 8'd192, 8'd138, 8'd143, 8'd93, 8'd137, 8'd90, 8'd92, 8'd92, 8'd154, 8'd129, 8'd110, 8'd148, 8'd178, 8'd143, 8'd97, 8'd108, 8'd161, 8'd84, 8'd132, 8'd88, 8'd69, 8'd121, 8'd146, 8'd102, 8'd171, 8'd86, 8'd144, 8'd167, 8'd124, 8'd139, 8'd87, 8'd171, 8'd127, 8'd84, 8'd152, 8'd171, 8'd155, 8'd158, 8'd134, 8'd97, 8'd122, 8'd186, 8'd148, 8'd159, 8'd72, 8'd104, 8'd127, 8'd124, 8'd54, 8'd126, 8'd63, 8'd151, 8'd103, 8'd101, 8'd85, 8'd109, 8'd131, 8'd89, 8'd141, 8'd81, 8'd145, 8'd175, 8'd75, 8'd128, 8'd100, 8'd95, 8'd85, 8'd97, 8'd100, 8'd86, 8'd143, 8'd125, 8'd119, 8'd154, 8'd66, 8'd115, 8'd55, 8'd127, 8'd92, 8'd141, 8'd51, 8'd78, 8'd68, 8'd49, 8'd114, 8'd74, 8'd149, 8'd72, 8'd145, 8'd118, 8'd71, 8'd101, 8'd139, 8'd94, 8'd120, 8'd150, 8'd105, 8'd121, 8'd117, 8'd116, 8'd163, 8'd141, 8'd130, 8'd77, 8'd100, 8'd96, 8'd80, 8'd93, 8'd122, 8'd135, 8'd84, 8'd87, 8'd62, 8'd106, 8'd143, 8'd81, 8'd119, 8'd96, 8'd134, 8'd145, 8'd149, 8'd127, 8'd75, 8'd143, 8'd122, 8'd144, 8'd112, 8'd139, 8'd161, 8'd131, 8'd115, 8'd139, 8'd141, 8'd70, 8'd69, 8'd62, 8'd101, 8'd29, 8'd121, 8'd40, 8'd97, 8'd84, 8'd138, 8'd63, 8'd135, 8'd117, 8'd55, 8'd131, 8'd97, 8'd85, 8'd164, 8'd78, 8'd83, 8'd151, 8'd163, 8'd159, 8'd124, 8'd112, 8'd94, 8'd149, 8'd123, 8'd125, 8'd153, 8'd143, 8'd117, 8'd110, 8'd121, 8'd83, 8'd79, 8'd151, 8'd112, 8'd164, 8'd156, 8'd97, 8'd167, 8'd82, 8'd93, 8'd141, 8'd86, 8'd156, 8'd175, 8'd95, 8'd141, 8'd112, 8'd110, 8'd154, 8'd140, 8'd156, 8'd91, 8'd159, 8'd169, 8'd119, 8'd144, 8'd160, 8'd100, 8'd119, 8'd116, 8'd172, 8'd84, 8'd154, 8'd132, 8'd139, 8'd85, 8'd149, 8'd144, 8'd184, 8'd148, 8'd91, 8'd158, 8'd117, 8'd70, 8'd140, 8'd158, 8'd80, 8'd87, 8'd134, 8'd96, 8'd71, 8'd102, 8'd134, 8'd98, 8'd95, 8'd111, 8'd88, 8'd133, 8'd127, 8'd110, 8'd105, 8'd144, 8'd118, 8'd78, 8'd118, 8'd131, 8'd79, 8'd140, 8'd77, 8'd141, 8'd125, 8'd73, 8'd158, 8'd73})
) cell_0_41 (
    .clk(clk),
    .input_index(index_0_40_41),
    .input_value(value_0_40_41),
    .input_result(result_0_40_41),
    .input_enable(enable_0_40_41),
    .output_index(index_0_41_42),
    .output_value(value_0_41_42),
    .output_result(result_0_41_42),
    .output_enable(enable_0_41_42)
);

wire [10-1:0] index_0_42_43;
wire [`DATA_WIDTH-1:0] value_0_42_43;
wire [`DATA_WIDTH*4:0] result_0_42_43;
wire enable_0_42_43;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd81, 8'd150, 8'd113, 8'd70, 8'd157, 8'd72, 8'd113, 8'd128, 8'd86, 8'd154, 8'd126, 8'd103, 8'd178, 8'd189, 8'd171, 8'd176, 8'd137, 8'd145, 8'd147, 8'd171, 8'd111, 8'd116, 8'd150, 8'd79, 8'd111, 8'd150, 8'd137, 8'd84, 8'd162, 8'd79, 8'd130, 8'd121, 8'd159, 8'd190, 8'd130, 8'd152, 8'd116, 8'd167, 8'd182, 8'd149, 8'd184, 8'd204, 8'd215, 8'd224, 8'd185, 8'd166, 8'd174, 8'd175, 8'd115, 8'd116, 8'd82, 8'd138, 8'd160, 8'd139, 8'd128, 8'd155, 8'd93, 8'd104, 8'd100, 8'd173, 8'd149, 8'd176, 8'd115, 8'd169, 8'd194, 8'd169, 8'd124, 8'd118, 8'd113, 8'd121, 8'd195, 8'd203, 8'd123, 8'd178, 8'd145, 8'd159, 8'd113, 8'd166, 8'd163, 8'd109, 8'd87, 8'd122, 8'd81, 8'd160, 8'd129, 8'd102, 8'd135, 8'd98, 8'd164, 8'd117, 8'd118, 8'd143, 8'd123, 8'd106, 8'd72, 8'd94, 8'd128, 8'd144, 8'd138, 8'd129, 8'd145, 8'd92, 8'd117, 8'd83, 8'd104, 8'd136, 8'd146, 8'd131, 8'd180, 8'd154, 8'd81, 8'd98, 8'd141, 8'd73, 8'd98, 8'd150, 8'd99, 8'd101, 8'd66, 8'd87, 8'd138, 8'd65, 8'd73, 8'd106, 8'd153, 8'd114, 8'd116, 8'd104, 8'd104, 8'd142, 8'd83, 8'd173, 8'd111, 8'd85, 8'd111, 8'd106, 8'd156, 8'd143, 8'd87, 8'd167, 8'd146, 8'd98, 8'd127, 8'd144, 8'd95, 8'd162, 8'd84, 8'd82, 8'd132, 8'd150, 8'd86, 8'd72, 8'd103, 8'd141, 8'd181, 8'd96, 8'd156, 8'd99, 8'd114, 8'd147, 8'd123, 8'd156, 8'd147, 8'd147, 8'd137, 8'd61, 8'd71, 8'd151, 8'd96, 8'd85, 8'd86, 8'd143, 8'd94, 8'd112, 8'd85, 8'd119, 8'd145, 8'd62, 8'd97, 8'd124, 8'd77, 8'd77, 8'd156, 8'd91, 8'd175, 8'd148, 8'd85, 8'd139, 8'd152, 8'd84, 8'd95, 8'd83, 8'd104, 8'd152, 8'd104, 8'd75, 8'd127, 8'd65, 8'd128, 8'd146, 8'd139, 8'd77, 8'd145, 8'd143, 8'd126, 8'd143, 8'd103, 8'd64, 8'd93, 8'd66, 8'd137, 8'd158, 8'd113, 8'd140, 8'd115, 8'd125, 8'd83, 8'd162, 8'd133, 8'd89, 8'd156, 8'd130, 8'd125, 8'd150, 8'd110, 8'd77, 8'd43, 8'd100, 8'd133, 8'd80, 8'd134, 8'd160, 8'd96, 8'd147, 8'd122, 8'd86, 8'd134, 8'd55, 8'd138, 8'd158, 8'd84, 8'd161, 8'd75, 8'd113, 8'd157, 8'd170, 8'd147, 8'd167, 8'd132, 8'd153, 8'd161, 8'd164, 8'd130, 8'd145, 8'd45, 8'd101, 8'd82, 8'd98, 8'd96, 8'd93, 8'd130, 8'd105, 8'd157, 8'd111, 8'd121, 8'd72, 8'd100, 8'd66, 8'd129, 8'd77, 8'd159, 8'd150, 8'd88, 8'd140, 8'd89, 8'd92, 8'd131, 8'd127, 8'd87, 8'd116, 8'd169, 8'd98, 8'd107, 8'd114, 8'd107, 8'd80, 8'd167, 8'd152, 8'd91, 8'd126, 8'd157, 8'd70, 8'd98, 8'd121, 8'd30, 8'd84, 8'd101, 8'd127, 8'd124, 8'd122, 8'd83, 8'd140, 8'd135, 8'd90, 8'd88, 8'd75, 8'd123, 8'd70, 8'd132, 8'd66, 8'd71, 8'd143, 8'd145, 8'd101, 8'd159, 8'd120, 8'd102, 8'd155, 8'd156, 8'd63, 8'd94, 8'd52, 8'd31, 8'd97, 8'd91, 8'd77, 8'd158, 8'd84, 8'd108, 8'd84, 8'd162, 8'd84, 8'd101, 8'd120, 8'd84, 8'd133, 8'd62, 8'd128, 8'd72, 8'd87, 8'd86, 8'd167, 8'd158, 8'd78, 8'd127, 8'd78, 8'd143, 8'd129, 8'd42, 8'd117, 8'd90, 8'd120, 8'd138, 8'd148, 8'd89, 8'd103, 8'd159, 8'd78, 8'd160, 8'd108, 8'd115, 8'd68, 8'd118, 8'd99, 8'd139, 8'd48, 8'd146, 8'd138, 8'd167, 8'd136, 8'd133, 8'd131, 8'd160, 8'd160, 8'd61, 8'd80, 8'd117, 8'd96, 8'd108, 8'd81, 8'd66, 8'd135, 8'd111, 8'd92, 8'd80, 8'd87, 8'd116, 8'd137, 8'd94, 8'd94, 8'd177, 8'd119, 8'd159, 8'd83, 8'd75, 8'd81, 8'd81, 8'd85, 8'd135, 8'd100, 8'd86, 8'd152, 8'd131, 8'd127, 8'd59, 8'd78, 8'd134, 8'd150, 8'd105, 8'd111, 8'd87, 8'd139, 8'd102, 8'd148, 8'd130, 8'd146, 8'd141, 8'd182, 8'd96, 8'd116, 8'd144, 8'd110, 8'd113, 8'd132, 8'd93, 8'd93, 8'd155, 8'd102, 8'd129, 8'd91, 8'd108, 8'd99, 8'd82, 8'd131, 8'd105, 8'd85, 8'd120, 8'd99, 8'd103, 8'd163, 8'd174, 8'd158, 8'd96, 8'd134, 8'd120, 8'd182, 8'd184, 8'd157, 8'd128, 8'd114, 8'd122, 8'd164, 8'd116, 8'd77, 8'd127, 8'd141, 8'd151, 8'd94, 8'd142, 8'd61, 8'd102, 8'd100, 8'd172, 8'd115, 8'd126, 8'd115, 8'd76, 8'd174, 8'd150, 8'd124, 8'd132, 8'd150, 8'd140, 8'd120, 8'd110, 8'd95, 8'd117, 8'd142, 8'd170, 8'd169, 8'd167, 8'd173, 8'd106, 8'd102, 8'd167, 8'd168, 8'd85, 8'd125, 8'd175, 8'd127, 8'd143, 8'd183, 8'd137, 8'd97, 8'd165, 8'd91, 8'd127, 8'd109, 8'd111, 8'd90, 8'd141, 8'd156, 8'd109, 8'd166, 8'd107, 8'd150, 8'd164, 8'd207, 8'd139, 8'd139, 8'd83, 8'd86, 8'd171, 8'd170, 8'd176, 8'd120, 8'd129, 8'd134, 8'd148, 8'd88, 8'd131, 8'd151, 8'd154, 8'd109, 8'd166, 8'd113, 8'd158, 8'd103, 8'd163, 8'd117, 8'd136, 8'd162, 8'd171, 8'd128, 8'd160, 8'd132, 8'd193, 8'd147, 8'd148, 8'd130, 8'd173, 8'd135, 8'd100, 8'd117, 8'd112, 8'd125, 8'd157, 8'd137, 8'd128, 8'd73, 8'd123, 8'd156, 8'd75, 8'd154, 8'd136, 8'd78, 8'd147, 8'd74, 8'd151, 8'd175, 8'd88, 8'd143, 8'd172, 8'd86, 8'd180, 8'd79, 8'd117, 8'd166, 8'd126, 8'd184, 8'd179, 8'd131, 8'd164, 8'd114, 8'd87, 8'd146, 8'd111, 8'd173, 8'd111, 8'd158, 8'd99, 8'd161, 8'd75, 8'd54, 8'd113, 8'd90, 8'd79, 8'd104, 8'd132, 8'd132, 8'd144, 8'd85, 8'd161, 8'd74, 8'd100, 8'd146, 8'd99, 8'd182, 8'd99, 8'd172, 8'd129, 8'd90, 8'd176, 8'd113, 8'd92, 8'd130, 8'd137, 8'd81, 8'd158, 8'd145, 8'd75, 8'd138, 8'd125, 8'd132, 8'd83, 8'd71, 8'd83, 8'd127, 8'd169, 8'd102, 8'd74, 8'd159, 8'd148, 8'd121, 8'd155, 8'd79, 8'd117, 8'd85, 8'd97, 8'd141, 8'd160, 8'd76, 8'd149, 8'd120, 8'd60, 8'd97, 8'd101, 8'd136, 8'd77, 8'd96, 8'd92, 8'd145, 8'd158, 8'd134, 8'd106, 8'd108, 8'd123, 8'd86, 8'd89, 8'd114, 8'd65, 8'd71, 8'd146, 8'd135, 8'd78, 8'd146, 8'd162, 8'd157, 8'd145, 8'd77, 8'd156, 8'd131, 8'd136, 8'd119, 8'd74, 8'd142, 8'd131, 8'd79, 8'd100, 8'd122, 8'd114, 8'd77, 8'd143, 8'd90, 8'd132, 8'd122, 8'd74, 8'd131, 8'd83, 8'd124, 8'd80, 8'd79, 8'd115, 8'd143, 8'd71, 8'd118, 8'd81, 8'd108, 8'd73, 8'd73, 8'd136, 8'd103, 8'd111, 8'd150, 8'd126, 8'd126, 8'd169, 8'd103, 8'd145, 8'd95, 8'd124, 8'd134, 8'd92, 8'd156, 8'd105, 8'd158, 8'd84, 8'd70, 8'd99, 8'd135, 8'd140, 8'd84, 8'd101, 8'd102, 8'd107, 8'd89, 8'd130, 8'd168, 8'd96, 8'd167, 8'd140, 8'd122, 8'd86, 8'd112, 8'd85, 8'd141, 8'd137, 8'd163, 8'd166, 8'd79, 8'd141, 8'd88, 8'd91, 8'd159, 8'd102, 8'd181, 8'd87, 8'd166, 8'd117, 8'd149, 8'd144, 8'd136, 8'd182, 8'd169, 8'd157, 8'd145, 8'd167, 8'd148, 8'd149, 8'd158, 8'd116, 8'd133, 8'd114, 8'd163, 8'd154, 8'd101, 8'd159, 8'd88, 8'd107, 8'd133, 8'd118, 8'd139, 8'd101, 8'd152, 8'd166, 8'd100, 8'd112, 8'd117, 8'd163, 8'd76, 8'd164, 8'd148, 8'd150, 8'd123, 8'd104, 8'd121, 8'd111, 8'd93, 8'd110, 8'd98, 8'd157, 8'd111, 8'd91, 8'd92})
) cell_0_42 (
    .clk(clk),
    .input_index(index_0_41_42),
    .input_value(value_0_41_42),
    .input_result(result_0_41_42),
    .input_enable(enable_0_41_42),
    .output_index(index_0_42_43),
    .output_value(value_0_42_43),
    .output_result(result_0_42_43),
    .output_enable(enable_0_42_43)
);

wire [10-1:0] index_0_43_44;
wire [`DATA_WIDTH-1:0] value_0_43_44;
wire [`DATA_WIDTH*4:0] result_0_43_44;
wire enable_0_43_44;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd125, 8'd107, 8'd155, 8'd169, 8'd170, 8'd124, 8'd175, 8'd100, 8'd91, 8'd180, 8'd186, 8'd106, 8'd181, 8'd111, 8'd119, 8'd164, 8'd96, 8'd101, 8'd125, 8'd161, 8'd130, 8'd145, 8'd150, 8'd138, 8'd111, 8'd122, 8'd102, 8'd103, 8'd78, 8'd138, 8'd156, 8'd102, 8'd150, 8'd141, 8'd88, 8'd62, 8'd55, 8'd108, 8'd131, 8'd125, 8'd94, 8'd101, 8'd124, 8'd72, 8'd94, 8'd81, 8'd57, 8'd96, 8'd62, 8'd110, 8'd62, 8'd147, 8'd71, 8'd108, 8'd162, 8'd96, 8'd121, 8'd96, 8'd150, 8'd114, 8'd77, 8'd62, 8'd42, 8'd125, 8'd97, 8'd126, 8'd108, 8'd62, 8'd127, 8'd82, 8'd79, 8'd112, 8'd96, 8'd69, 8'd65, 8'd62, 8'd118, 8'd69, 8'd120, 8'd99, 8'd67, 8'd135, 8'd97, 8'd91, 8'd167, 8'd174, 8'd106, 8'd99, 8'd71, 8'd141, 8'd126, 8'd97, 8'd127, 8'd161, 8'd125, 8'd79, 8'd142, 8'd116, 8'd81, 8'd157, 8'd152, 8'd116, 8'd80, 8'd68, 8'd86, 8'd77, 8'd83, 8'd90, 8'd90, 8'd97, 8'd135, 8'd118, 8'd92, 8'd94, 8'd91, 8'd117, 8'd73, 8'd143, 8'd160, 8'd167, 8'd156, 8'd121, 8'd166, 8'd115, 8'd164, 8'd121, 8'd104, 8'd81, 8'd120, 8'd97, 8'd117, 8'd146, 8'd81, 8'd90, 8'd151, 8'd147, 8'd131, 8'd73, 8'd80, 8'd153, 8'd78, 8'd124, 8'd113, 8'd181, 8'd173, 8'd169, 8'd156, 8'd148, 8'd151, 8'd124, 8'd82, 8'd93, 8'd96, 8'd142, 8'd112, 8'd80, 8'd108, 8'd77, 8'd147, 8'd92, 8'd86, 8'd111, 8'd77, 8'd94, 8'd104, 8'd146, 8'd100, 8'd155, 8'd73, 8'd109, 8'd143, 8'd128, 8'd129, 8'd106, 8'd166, 8'd83, 8'd120, 8'd118, 8'd81, 8'd143, 8'd141, 8'd106, 8'd136, 8'd170, 8'd151, 8'd149, 8'd179, 8'd106, 8'd155, 8'd137, 8'd105, 8'd144, 8'd129, 8'd134, 8'd142, 8'd94, 8'd131, 8'd134, 8'd109, 8'd141, 8'd163, 8'd124, 8'd168, 8'd110, 8'd93, 8'd145, 8'd119, 8'd162, 8'd93, 8'd121, 8'd88, 8'd107, 8'd105, 8'd120, 8'd116, 8'd158, 8'd141, 8'd98, 8'd151, 8'd137, 8'd162, 8'd171, 8'd111, 8'd78, 8'd106, 8'd198, 8'd131, 8'd163, 8'd118, 8'd171, 8'd105, 8'd154, 8'd96, 8'd106, 8'd97, 8'd163, 8'd142, 8'd171, 8'd110, 8'd105, 8'd126, 8'd124, 8'd93, 8'd73, 8'd112, 8'd127, 8'd156, 8'd166, 8'd116, 8'd148, 8'd119, 8'd78, 8'd130, 8'd132, 8'd179, 8'd117, 8'd125, 8'd125, 8'd158, 8'd112, 8'd109, 8'd126, 8'd103, 8'd126, 8'd118, 8'd124, 8'd180, 8'd157, 8'd94, 8'd116, 8'd99, 8'd125, 8'd109, 8'd123, 8'd113, 8'd111, 8'd152, 8'd125, 8'd76, 8'd148, 8'd112, 8'd114, 8'd128, 8'd135, 8'd150, 8'd162, 8'd109, 8'd127, 8'd85, 8'd79, 8'd81, 8'd154, 8'd162, 8'd154, 8'd160, 8'd109, 8'd102, 8'd152, 8'd151, 8'd151, 8'd103, 8'd87, 8'd139, 8'd79, 8'd170, 8'd149, 8'd115, 8'd121, 8'd160, 8'd122, 8'd186, 8'd91, 8'd74, 8'd86, 8'd125, 8'd75, 8'd127, 8'd152, 8'd91, 8'd159, 8'd133, 8'd194, 8'd185, 8'd193, 8'd90, 8'd107, 8'd131, 8'd115, 8'd134, 8'd85, 8'd78, 8'd174, 8'd107, 8'd141, 8'd119, 8'd149, 8'd136, 8'd190, 8'd129, 8'd161, 8'd60, 8'd114, 8'd127, 8'd101, 8'd128, 8'd146, 8'd152, 8'd148, 8'd134, 8'd119, 8'd160, 8'd94, 8'd102, 8'd60, 8'd157, 8'd160, 8'd118, 8'd109, 8'd78, 8'd148, 8'd151, 8'd81, 8'd118, 8'd112, 8'd96, 8'd164, 8'd147, 8'd171, 8'd111, 8'd82, 8'd118, 8'd86, 8'd181, 8'd113, 8'd117, 8'd122, 8'd81, 8'd160, 8'd100, 8'd69, 8'd127, 8'd89, 8'd101, 8'd107, 8'd145, 8'd72, 8'd119, 8'd126, 8'd110, 8'd184, 8'd159, 8'd138, 8'd179, 8'd168, 8'd162, 8'd108, 8'd118, 8'd130, 8'd102, 8'd97, 8'd124, 8'd130, 8'd132, 8'd146, 8'd86, 8'd147, 8'd89, 8'd80, 8'd112, 8'd94, 8'd85, 8'd67, 8'd75, 8'd96, 8'd107, 8'd111, 8'd112, 8'd95, 8'd164, 8'd98, 8'd85, 8'd124, 8'd183, 8'd172, 8'd90, 8'd84, 8'd107, 8'd96, 8'd76, 8'd90, 8'd150, 8'd134, 8'd101, 8'd73, 8'd59, 8'd47, 8'd76, 8'd68, 8'd124, 8'd107, 8'd53, 8'd99, 8'd112, 8'd62, 8'd95, 8'd90, 8'd137, 8'd106, 8'd144, 8'd103, 8'd116, 8'd118, 8'd63, 8'd93, 8'd156, 8'd123, 8'd123, 8'd100, 8'd115, 8'd118, 8'd79, 8'd99, 8'd33, 8'd42, 8'd141, 8'd93, 8'd96, 8'd91, 8'd78, 8'd101, 8'd161, 8'd111, 8'd139, 8'd106, 8'd152, 8'd171, 8'd88, 8'd96, 8'd36, 8'd35, 8'd121, 8'd105, 8'd161, 8'd94, 8'd148, 8'd94, 8'd138, 8'd125, 8'd88, 8'd73, 8'd78, 8'd110, 8'd115, 8'd74, 8'd155, 8'd73, 8'd157, 8'd136, 8'd159, 8'd151, 8'd100, 8'd100, 8'd139, 8'd148, 8'd136, 8'd97, 8'd40, 8'd21, 8'd140, 8'd161, 8'd126, 8'd84, 8'd90, 8'd123, 8'd128, 8'd94, 8'd145, 8'd72, 8'd141, 8'd158, 8'd117, 8'd103, 8'd100, 8'd95, 8'd169, 8'd137, 8'd133, 8'd115, 8'd176, 8'd128, 8'd143, 8'd135, 8'd140, 8'd133, 8'd126, 8'd96, 8'd144, 8'd124, 8'd107, 8'd119, 8'd152, 8'd157, 8'd77, 8'd140, 8'd69, 8'd134, 8'd154, 8'd107, 8'd104, 8'd167, 8'd115, 8'd145, 8'd91, 8'd173, 8'd192, 8'd132, 8'd165, 8'd133, 8'd113, 8'd108, 8'd124, 8'd125, 8'd76, 8'd65, 8'd153, 8'd89, 8'd109, 8'd74, 8'd75, 8'd131, 8'd53, 8'd138, 8'd142, 8'd78, 8'd73, 8'd150, 8'd140, 8'd155, 8'd182, 8'd141, 8'd135, 8'd185, 8'd162, 8'd153, 8'd157, 8'd141, 8'd159, 8'd125, 8'd103, 8'd126, 8'd157, 8'd75, 8'd98, 8'd74, 8'd87, 8'd104, 8'd82, 8'd102, 8'd91, 8'd133, 8'd144, 8'd114, 8'd124, 8'd156, 8'd115, 8'd137, 8'd106, 8'd103, 8'd148, 8'd130, 8'd92, 8'd111, 8'd165, 8'd129, 8'd149, 8'd131, 8'd105, 8'd84, 8'd133, 8'd62, 8'd95, 8'd109, 8'd106, 8'd152, 8'd107, 8'd161, 8'd91, 8'd116, 8'd108, 8'd103, 8'd85, 8'd106, 8'd93, 8'd176, 8'd95, 8'd104, 8'd152, 8'd115, 8'd188, 8'd116, 8'd128, 8'd73, 8'd167, 8'd125, 8'd154, 8'd144, 8'd154, 8'd122, 8'd50, 8'd108, 8'd155, 8'd120, 8'd111, 8'd165, 8'd103, 8'd124, 8'd98, 8'd173, 8'd90, 8'd128, 8'd135, 8'd137, 8'd150, 8'd113, 8'd107, 8'd87, 8'd178, 8'd85, 8'd100, 8'd91, 8'd123, 8'd127, 8'd129, 8'd135, 8'd125, 8'd134, 8'd134, 8'd97, 8'd76, 8'd129, 8'd127, 8'd104, 8'd128, 8'd82, 8'd96, 8'd115, 8'd104, 8'd149, 8'd136, 8'd105, 8'd170, 8'd84, 8'd64, 8'd68, 8'd94, 8'd82, 8'd81, 8'd133, 8'd152, 8'd113, 8'd167, 8'd95, 8'd108, 8'd167, 8'd94, 8'd98, 8'd81, 8'd64, 8'd88, 8'd57, 8'd151, 8'd172, 8'd101, 8'd122, 8'd147, 8'd85, 8'd111, 8'd128, 8'd146, 8'd90, 8'd53, 8'd108, 8'd91, 8'd154, 8'd161, 8'd86, 8'd102, 8'd99, 8'd100, 8'd130, 8'd101, 8'd155, 8'd144, 8'd68, 8'd112, 8'd89, 8'd74, 8'd108, 8'd137, 8'd89, 8'd118, 8'd83, 8'd94, 8'd95, 8'd114, 8'd111, 8'd59, 8'd59, 8'd93, 8'd121, 8'd90, 8'd140, 8'd120, 8'd142, 8'd85, 8'd120, 8'd98, 8'd73, 8'd132, 8'd82, 8'd92, 8'd112, 8'd113, 8'd156, 8'd87, 8'd75, 8'd113, 8'd129, 8'd113, 8'd88, 8'd72, 8'd97, 8'd147, 8'd97, 8'd149, 8'd127, 8'd155, 8'd147, 8'd147, 8'd87, 8'd112, 8'd146, 8'd148, 8'd123})
) cell_0_43 (
    .clk(clk),
    .input_index(index_0_42_43),
    .input_value(value_0_42_43),
    .input_result(result_0_42_43),
    .input_enable(enable_0_42_43),
    .output_index(index_0_43_44),
    .output_value(value_0_43_44),
    .output_result(result_0_43_44),
    .output_enable(enable_0_43_44)
);

wire [10-1:0] index_0_44_45;
wire [`DATA_WIDTH-1:0] value_0_44_45;
wire [`DATA_WIDTH*4:0] result_0_44_45;
wire enable_0_44_45;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd81, 8'd155, 8'd159, 8'd123, 8'd105, 8'd135, 8'd116, 8'd150, 8'd164, 8'd179, 8'd164, 8'd177, 8'd182, 8'd193, 8'd164, 8'd146, 8'd171, 8'd175, 8'd154, 8'd128, 8'd151, 8'd163, 8'd134, 8'd159, 8'd71, 8'd76, 8'd123, 8'd160, 8'd135, 8'd99, 8'd168, 8'd81, 8'd117, 8'd169, 8'd74, 8'd77, 8'd180, 8'd115, 8'd191, 8'd154, 8'd147, 8'd131, 8'd191, 8'd137, 8'd131, 8'd95, 8'd99, 8'd127, 8'd174, 8'd107, 8'd142, 8'd102, 8'd121, 8'd113, 8'd124, 8'd112, 8'd136, 8'd92, 8'd137, 8'd66, 8'd93, 8'd122, 8'd135, 8'd111, 8'd113, 8'd139, 8'd139, 8'd109, 8'd126, 8'd96, 8'd124, 8'd89, 8'd82, 8'd70, 8'd61, 8'd68, 8'd94, 8'd100, 8'd55, 8'd132, 8'd73, 8'd161, 8'd151, 8'd85, 8'd134, 8'd76, 8'd84, 8'd151, 8'd72, 8'd90, 8'd105, 8'd73, 8'd122, 8'd149, 8'd111, 8'd155, 8'd105, 8'd132, 8'd149, 8'd94, 8'd159, 8'd116, 8'd126, 8'd139, 8'd65, 8'd79, 8'd122, 8'd126, 8'd106, 8'd82, 8'd100, 8'd102, 8'd83, 8'd64, 8'd70, 8'd111, 8'd67, 8'd128, 8'd102, 8'd155, 8'd109, 8'd131, 8'd131, 8'd156, 8'd145, 8'd153, 8'd151, 8'd89, 8'd157, 8'd67, 8'd110, 8'd112, 8'd160, 8'd88, 8'd64, 8'd129, 8'd126, 8'd96, 8'd84, 8'd115, 8'd90, 8'd93, 8'd78, 8'd77, 8'd118, 8'd107, 8'd116, 8'd103, 8'd153, 8'd127, 8'd162, 8'd168, 8'd113, 8'd100, 8'd93, 8'd142, 8'd125, 8'd81, 8'd163, 8'd139, 8'd75, 8'd121, 8'd151, 8'd78, 8'd106, 8'd153, 8'd147, 8'd124, 8'd107, 8'd152, 8'd128, 8'd142, 8'd78, 8'd91, 8'd138, 8'd134, 8'd111, 8'd104, 8'd139, 8'd92, 8'd78, 8'd147, 8'd174, 8'd160, 8'd148, 8'd119, 8'd96, 8'd99, 8'd93, 8'd83, 8'd110, 8'd83, 8'd65, 8'd53, 8'd150, 8'd145, 8'd123, 8'd106, 8'd146, 8'd101, 8'd166, 8'd124, 8'd129, 8'd159, 8'd171, 8'd111, 8'd75, 8'd131, 8'd139, 8'd160, 8'd106, 8'd142, 8'd117, 8'd132, 8'd148, 8'd171, 8'd172, 8'd67, 8'd86, 8'd61, 8'd121, 8'd72, 8'd161, 8'd112, 8'd95, 8'd131, 8'd134, 8'd102, 8'd134, 8'd109, 8'd127, 8'd139, 8'd172, 8'd130, 8'd103, 8'd132, 8'd134, 8'd99, 8'd120, 8'd148, 8'd125, 8'd183, 8'd118, 8'd80, 8'd90, 8'd152, 8'd80, 8'd121, 8'd43, 8'd119, 8'd84, 8'd152, 8'd140, 8'd133, 8'd76, 8'd140, 8'd139, 8'd112, 8'd73, 8'd74, 8'd134, 8'd149, 8'd82, 8'd77, 8'd113, 8'd126, 8'd116, 8'd124, 8'd191, 8'd159, 8'd104, 8'd152, 8'd79, 8'd143, 8'd66, 8'd61, 8'd98, 8'd118, 8'd161, 8'd115, 8'd137, 8'd138, 8'd112, 8'd148, 8'd98, 8'd105, 8'd82, 8'd86, 8'd140, 8'd118, 8'd106, 8'd96, 8'd97, 8'd115, 8'd175, 8'd105, 8'd202, 8'd136, 8'd164, 8'd142, 8'd88, 8'd96, 8'd154, 8'd67, 8'd83, 8'd140, 8'd151, 8'd84, 8'd96, 8'd93, 8'd152, 8'd102, 8'd139, 8'd71, 8'd127, 8'd62, 8'd85, 8'd124, 8'd152, 8'd148, 8'd78, 8'd95, 8'd90, 8'd111, 8'd182, 8'd149, 8'd90, 8'd152, 8'd176, 8'd118, 8'd158, 8'd132, 8'd125, 8'd143, 8'd120, 8'd96, 8'd63, 8'd120, 8'd127, 8'd83, 8'd110, 8'd161, 8'd128, 8'd96, 8'd59, 8'd95, 8'd63, 8'd156, 8'd126, 8'd134, 8'd92, 8'd133, 8'd119, 8'd72, 8'd106, 8'd158, 8'd148, 8'd97, 8'd136, 8'd122, 8'd94, 8'd87, 8'd150, 8'd118, 8'd64, 8'd53, 8'd143, 8'd175, 8'd175, 8'd123, 8'd169, 8'd86, 8'd142, 8'd100, 8'd109, 8'd117, 8'd135, 8'd125, 8'd87, 8'd155, 8'd150, 8'd102, 8'd82, 8'd69, 8'd83, 8'd150, 8'd96, 8'd131, 8'd128, 8'd174, 8'd138, 8'd83, 8'd66, 8'd51, 8'd109, 8'd142, 8'd142, 8'd120, 8'd142, 8'd168, 8'd156, 8'd114, 8'd151, 8'd66, 8'd147, 8'd113, 8'd105, 8'd114, 8'd136, 8'd57, 8'd159, 8'd138, 8'd147, 8'd132, 8'd121, 8'd133, 8'd147, 8'd103, 8'd119, 8'd110, 8'd76, 8'd127, 8'd85, 8'd137, 8'd207, 8'd171, 8'd120, 8'd162, 8'd138, 8'd93, 8'd110, 8'd155, 8'd55, 8'd87, 8'd148, 8'd138, 8'd160, 8'd151, 8'd117, 8'd121, 8'd139, 8'd120, 8'd163, 8'd86, 8'd138, 8'd114, 8'd88, 8'd86, 8'd136, 8'd53, 8'd88, 8'd141, 8'd118, 8'd144, 8'd99, 8'd158, 8'd167, 8'd83, 8'd71, 8'd76, 8'd58, 8'd85, 8'd94, 8'd97, 8'd86, 8'd150, 8'd157, 8'd167, 8'd154, 8'd87, 8'd145, 8'd152, 8'd68, 8'd179, 8'd108, 8'd147, 8'd142, 8'd116, 8'd116, 8'd113, 8'd143, 8'd114, 8'd102, 8'd126, 8'd138, 8'd85, 8'd153, 8'd56, 8'd139, 8'd148, 8'd81, 8'd104, 8'd119, 8'd99, 8'd94, 8'd92, 8'd112, 8'd89, 8'd85, 8'd123, 8'd77, 8'd79, 8'd155, 8'd85, 8'd112, 8'd122, 8'd65, 8'd71, 8'd100, 8'd153, 8'd141, 8'd158, 8'd88, 8'd85, 8'd108, 8'd108, 8'd73, 8'd91, 8'd84, 8'd90, 8'd82, 8'd153, 8'd128, 8'd109, 8'd175, 8'd139, 8'd91, 8'd157, 8'd100, 8'd145, 8'd129, 8'd164, 8'd129, 8'd81, 8'd135, 8'd78, 8'd145, 8'd124, 8'd79, 8'd88, 8'd144, 8'd69, 8'd89, 8'd159, 8'd89, 8'd73, 8'd132, 8'd130, 8'd86, 8'd100, 8'd147, 8'd160, 8'd176, 8'd124, 8'd145, 8'd111, 8'd140, 8'd107, 8'd75, 8'd155, 8'd86, 8'd78, 8'd102, 8'd144, 8'd132, 8'd87, 8'd97, 8'd82, 8'd119, 8'd84, 8'd74, 8'd137, 8'd70, 8'd145, 8'd89, 8'd102, 8'd112, 8'd145, 8'd143, 8'd128, 8'd96, 8'd89, 8'd153, 8'd138, 8'd145, 8'd92, 8'd128, 8'd155, 8'd135, 8'd102, 8'd162, 8'd127, 8'd83, 8'd168, 8'd109, 8'd148, 8'd147, 8'd140, 8'd99, 8'd117, 8'd97, 8'd103, 8'd137, 8'd149, 8'd134, 8'd100, 8'd148, 8'd139, 8'd111, 8'd139, 8'd126, 8'd137, 8'd86, 8'd116, 8'd114, 8'd94, 8'd71, 8'd106, 8'd151, 8'd159, 8'd133, 8'd97, 8'd172, 8'd114, 8'd142, 8'd139, 8'd83, 8'd144, 8'd121, 8'd145, 8'd137, 8'd137, 8'd96, 8'd87, 8'd150, 8'd121, 8'd77, 8'd86, 8'd49, 8'd91, 8'd83, 8'd98, 8'd95, 8'd98, 8'd158, 8'd97, 8'd111, 8'd132, 8'd128, 8'd110, 8'd115, 8'd137, 8'd90, 8'd142, 8'd174, 8'd91, 8'd101, 8'd121, 8'd139, 8'd63, 8'd138, 8'd101, 8'd121, 8'd76, 8'd103, 8'd124, 8'd89, 8'd140, 8'd112, 8'd151, 8'd72, 8'd111, 8'd138, 8'd151, 8'd117, 8'd95, 8'd173, 8'd130, 8'd84, 8'd99, 8'd156, 8'd159, 8'd121, 8'd124, 8'd91, 8'd148, 8'd172, 8'd162, 8'd173, 8'd94, 8'd165, 8'd164, 8'd99, 8'd90, 8'd116, 8'd81, 8'd112, 8'd123, 8'd77, 8'd160, 8'd161, 8'd87, 8'd112, 8'd82, 8'd116, 8'd121, 8'd116, 8'd189, 8'd187, 8'd94, 8'd170, 8'd123, 8'd111, 8'd140, 8'd202, 8'd209, 8'd122, 8'd206, 8'd182, 8'd112, 8'd120, 8'd130, 8'd80, 8'd110, 8'd176, 8'd162, 8'd82, 8'd154, 8'd151, 8'd94, 8'd121, 8'd169, 8'd91, 8'd105, 8'd171, 8'd90, 8'd122, 8'd95, 8'd96, 8'd105, 8'd165, 8'd162, 8'd103, 8'd175, 8'd179, 8'd120, 8'd112, 8'd164, 8'd176, 8'd182, 8'd139, 8'd134, 8'd154, 8'd140, 8'd99, 8'd99, 8'd133, 8'd89, 8'd117, 8'd159, 8'd160, 8'd149, 8'd154, 8'd164, 8'd70, 8'd80, 8'd152, 8'd100, 8'd105, 8'd132, 8'd138, 8'd127, 8'd149, 8'd72, 8'd161, 8'd157, 8'd164, 8'd86, 8'd86, 8'd84, 8'd168, 8'd74, 8'd142, 8'd112})
) cell_0_44 (
    .clk(clk),
    .input_index(index_0_43_44),
    .input_value(value_0_43_44),
    .input_result(result_0_43_44),
    .input_enable(enable_0_43_44),
    .output_index(index_0_44_45),
    .output_value(value_0_44_45),
    .output_result(result_0_44_45),
    .output_enable(enable_0_44_45)
);

wire [10-1:0] index_0_45_46;
wire [`DATA_WIDTH-1:0] value_0_45_46;
wire [`DATA_WIDTH*4:0] result_0_45_46;
wire enable_0_45_46;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd135, 8'd99, 8'd80, 8'd97, 8'd89, 8'd100, 8'd152, 8'd116, 8'd136, 8'd117, 8'd177, 8'd136, 8'd121, 8'd197, 8'd187, 8'd180, 8'd120, 8'd173, 8'd83, 8'd152, 8'd114, 8'd143, 8'd88, 8'd113, 8'd87, 8'd71, 8'd156, 8'd111, 8'd148, 8'd122, 8'd168, 8'd117, 8'd153, 8'd85, 8'd158, 8'd132, 8'd99, 8'd101, 8'd138, 8'd135, 8'd182, 8'd144, 8'd109, 8'd157, 8'd148, 8'd178, 8'd166, 8'd163, 8'd141, 8'd123, 8'd133, 8'd64, 8'd124, 8'd146, 8'd79, 8'd102, 8'd169, 8'd166, 8'd87, 8'd166, 8'd116, 8'd113, 8'd73, 8'd93, 8'd163, 8'd125, 8'd148, 8'd162, 8'd125, 8'd147, 8'd94, 8'd119, 8'd134, 8'd168, 8'd170, 8'd111, 8'd126, 8'd157, 8'd129, 8'd120, 8'd112, 8'd60, 8'd138, 8'd99, 8'd158, 8'd141, 8'd128, 8'd141, 8'd97, 8'd80, 8'd60, 8'd138, 8'd120, 8'd122, 8'd135, 8'd171, 8'd109, 8'd185, 8'd194, 8'd128, 8'd180, 8'd119, 8'd82, 8'd151, 8'd78, 8'd110, 8'd109, 8'd92, 8'd129, 8'd116, 8'd165, 8'd137, 8'd138, 8'd96, 8'd167, 8'd175, 8'd93, 8'd159, 8'd102, 8'd100, 8'd68, 8'd147, 8'd86, 8'd100, 8'd119, 8'd149, 8'd141, 8'd117, 8'd135, 8'd107, 8'd123, 8'd93, 8'd109, 8'd97, 8'd87, 8'd83, 8'd124, 8'd139, 8'd113, 8'd162, 8'd133, 8'd83, 8'd90, 8'd139, 8'd191, 8'd133, 8'd76, 8'd76, 8'd90, 8'd102, 8'd133, 8'd69, 8'd141, 8'd91, 8'd110, 8'd181, 8'd132, 8'd156, 8'd180, 8'd173, 8'd83, 8'd89, 8'd122, 8'd88, 8'd63, 8'd91, 8'd132, 8'd83, 8'd156, 8'd176, 8'd106, 8'd95, 8'd193, 8'd141, 8'd172, 8'd129, 8'd85, 8'd109, 8'd58, 8'd88, 8'd65, 8'd165, 8'd174, 8'd98, 8'd97, 8'd84, 8'd108, 8'd174, 8'd145, 8'd100, 8'd91, 8'd152, 8'd123, 8'd70, 8'd109, 8'd136, 8'd127, 8'd88, 8'd126, 8'd92, 8'd142, 8'd161, 8'd145, 8'd148, 8'd85, 8'd87, 8'd70, 8'd136, 8'd92, 8'd122, 8'd156, 8'd176, 8'd161, 8'd92, 8'd168, 8'd168, 8'd106, 8'd95, 8'd163, 8'd106, 8'd142, 8'd133, 8'd82, 8'd78, 8'd96, 8'd97, 8'd139, 8'd164, 8'd93, 8'd177, 8'd145, 8'd138, 8'd87, 8'd103, 8'd135, 8'd106, 8'd140, 8'd104, 8'd96, 8'd141, 8'd119, 8'd121, 8'd171, 8'd131, 8'd126, 8'd89, 8'd114, 8'd138, 8'd82, 8'd165, 8'd157, 8'd151, 8'd151, 8'd155, 8'd189, 8'd119, 8'd172, 8'd163, 8'd86, 8'd130, 8'd133, 8'd63, 8'd159, 8'd116, 8'd160, 8'd81, 8'd78, 8'd116, 8'd137, 8'd129, 8'd173, 8'd123, 8'd133, 8'd149, 8'd185, 8'd160, 8'd73, 8'd69, 8'd120, 8'd84, 8'd164, 8'd190, 8'd148, 8'd179, 8'd124, 8'd96, 8'd127, 8'd112, 8'd108, 8'd144, 8'd123, 8'd177, 8'd85, 8'd118, 8'd115, 8'd108, 8'd104, 8'd103, 8'd83, 8'd107, 8'd96, 8'd146, 8'd184, 8'd153, 8'd83, 8'd141, 8'd145, 8'd93, 8'd140, 8'd191, 8'd179, 8'd164, 8'd175, 8'd112, 8'd134, 8'd132, 8'd161, 8'd132, 8'd107, 8'd90, 8'd129, 8'd36, 8'd135, 8'd97, 8'd100, 8'd108, 8'd113, 8'd171, 8'd172, 8'd173, 8'd146, 8'd134, 8'd83, 8'd128, 8'd82, 8'd145, 8'd136, 8'd141, 8'd127, 8'd130, 8'd156, 8'd108, 8'd100, 8'd100, 8'd148, 8'd130, 8'd99, 8'd89, 8'd42, 8'd102, 8'd79, 8'd123, 8'd65, 8'd151, 8'd169, 8'd126, 8'd95, 8'd168, 8'd123, 8'd154, 8'd124, 8'd102, 8'd143, 8'd157, 8'd95, 8'd146, 8'd111, 8'd166, 8'd159, 8'd165, 8'd75, 8'd165, 8'd160, 8'd107, 8'd93, 8'd79, 8'd109, 8'd32, 8'd91, 8'd64, 8'd79, 8'd154, 8'd98, 8'd160, 8'd146, 8'd68, 8'd80, 8'd99, 8'd153, 8'd137, 8'd162, 8'd123, 8'd89, 8'd113, 8'd166, 8'd147, 8'd93, 8'd148, 8'd107, 8'd83, 8'd89, 8'd117, 8'd119, 8'd48, 8'd98, 8'd73, 8'd68, 8'd120, 8'd106, 8'd154, 8'd92, 8'd113, 8'd136, 8'd110, 8'd105, 8'd103, 8'd147, 8'd183, 8'd110, 8'd127, 8'd82, 8'd125, 8'd162, 8'd122, 8'd150, 8'd156, 8'd151, 8'd154, 8'd144, 8'd141, 8'd156, 8'd85, 8'd124, 8'd110, 8'd131, 8'd92, 8'd140, 8'd81, 8'd86, 8'd149, 8'd110, 8'd108, 8'd100, 8'd155, 8'd165, 8'd180, 8'd110, 8'd143, 8'd139, 8'd153, 8'd136, 8'd154, 8'd154, 8'd86, 8'd89, 8'd170, 8'd183, 8'd124, 8'd131, 8'd61, 8'd53, 8'd64, 8'd111, 8'd123, 8'd168, 8'd89, 8'd81, 8'd132, 8'd160, 8'd104, 8'd173, 8'd137, 8'd157, 8'd161, 8'd119, 8'd78, 8'd134, 8'd161, 8'd163, 8'd193, 8'd189, 8'd140, 8'd103, 8'd113, 8'd155, 8'd177, 8'd133, 8'd118, 8'd136, 8'd101, 8'd166, 8'd178, 8'd129, 8'd147, 8'd183, 8'd100, 8'd156, 8'd96, 8'd147, 8'd147, 8'd162, 8'd187, 8'd154, 8'd144, 8'd93, 8'd138, 8'd217, 8'd185, 8'd213, 8'd130, 8'd142, 8'd192, 8'd161, 8'd162, 8'd103, 8'd89, 8'd79, 8'd166, 8'd159, 8'd166, 8'd147, 8'd165, 8'd120, 8'd192, 8'd85, 8'd177, 8'd115, 8'd147, 8'd172, 8'd131, 8'd165, 8'd136, 8'd96, 8'd83, 8'd151, 8'd141, 8'd142, 8'd140, 8'd126, 8'd185, 8'd118, 8'd170, 8'd157, 8'd101, 8'd120, 8'd130, 8'd169, 8'd103, 8'd200, 8'd168, 8'd140, 8'd179, 8'd142, 8'd105, 8'd137, 8'd107, 8'd153, 8'd124, 8'd102, 8'd168, 8'd92, 8'd68, 8'd100, 8'd157, 8'd152, 8'd102, 8'd166, 8'd133, 8'd135, 8'd126, 8'd168, 8'd100, 8'd83, 8'd94, 8'd141, 8'd91, 8'd191, 8'd104, 8'd140, 8'd134, 8'd141, 8'd118, 8'd80, 8'd137, 8'd165, 8'd152, 8'd121, 8'd107, 8'd81, 8'd82, 8'd130, 8'd116, 8'd81, 8'd116, 8'd173, 8'd92, 8'd104, 8'd142, 8'd113, 8'd86, 8'd87, 8'd172, 8'd89, 8'd90, 8'd169, 8'd178, 8'd107, 8'd147, 8'd83, 8'd88, 8'd147, 8'd67, 8'd103, 8'd90, 8'd97, 8'd75, 8'd104, 8'd175, 8'd180, 8'd156, 8'd66, 8'd138, 8'd154, 8'd80, 8'd73, 8'd91, 8'd123, 8'd134, 8'd161, 8'd90, 8'd170, 8'd95, 8'd128, 8'd104, 8'd135, 8'd143, 8'd120, 8'd140, 8'd138, 8'd56, 8'd74, 8'd121, 8'd98, 8'd157, 8'd135, 8'd153, 8'd171, 8'd77, 8'd122, 8'd60, 8'd135, 8'd123, 8'd117, 8'd76, 8'd99, 8'd101, 8'd115, 8'd156, 8'd116, 8'd111, 8'd108, 8'd137, 8'd105, 8'd127, 8'd72, 8'd126, 8'd49, 8'd58, 8'd159, 8'd145, 8'd146, 8'd109, 8'd116, 8'd170, 8'd132, 8'd105, 8'd52, 8'd137, 8'd140, 8'd128, 8'd147, 8'd122, 8'd70, 8'd50, 8'd71, 8'd64, 8'd152, 8'd129, 8'd93, 8'd139, 8'd149, 8'd95, 8'd96, 8'd96, 8'd99, 8'd84, 8'd138, 8'd122, 8'd80, 8'd77, 8'd96, 8'd167, 8'd79, 8'd140, 8'd83, 8'd115, 8'd121, 8'd43, 8'd52, 8'd121, 8'd99, 8'd125, 8'd132, 8'd88, 8'd102, 8'd139, 8'd56, 8'd53, 8'd146, 8'd153, 8'd152, 8'd65, 8'd159, 8'd83, 8'd133, 8'd130, 8'd148, 8'd145, 8'd155, 8'd99, 8'd74, 8'd94, 8'd101, 8'd152, 8'd54, 8'd69, 8'd102, 8'd88, 8'd119, 8'd93, 8'd144, 8'd83, 8'd95, 8'd99, 8'd136, 8'd54, 8'd105, 8'd124, 8'd90, 8'd100, 8'd76, 8'd83, 8'd118, 8'd169, 8'd77, 8'd96, 8'd91, 8'd158, 8'd152, 8'd165, 8'd115, 8'd152, 8'd142, 8'd101, 8'd134, 8'd127, 8'd115, 8'd78, 8'd146, 8'd74, 8'd142, 8'd147, 8'd137, 8'd111, 8'd105, 8'd136, 8'd152, 8'd149, 8'd132, 8'd154, 8'd107, 8'd110, 8'd72, 8'd75})
) cell_0_45 (
    .clk(clk),
    .input_index(index_0_44_45),
    .input_value(value_0_44_45),
    .input_result(result_0_44_45),
    .input_enable(enable_0_44_45),
    .output_index(index_0_45_46),
    .output_value(value_0_45_46),
    .output_result(result_0_45_46),
    .output_enable(enable_0_45_46)
);

wire [10-1:0] index_0_46_47;
wire [`DATA_WIDTH-1:0] value_0_46_47;
wire [`DATA_WIDTH*4:0] result_0_46_47;
wire enable_0_46_47;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd166, 8'd153, 8'd142, 8'd161, 8'd128, 8'd101, 8'd95, 8'd101, 8'd79, 8'd63, 8'd72, 8'd133, 8'd107, 8'd134, 8'd129, 8'd78, 8'd145, 8'd76, 8'd109, 8'd141, 8'd127, 8'd154, 8'd81, 8'd77, 8'd131, 8'd128, 8'd142, 8'd70, 8'd141, 8'd122, 8'd92, 8'd131, 8'd122, 8'd137, 8'd134, 8'd94, 8'd132, 8'd97, 8'd140, 8'd90, 8'd125, 8'd109, 8'd133, 8'd114, 8'd95, 8'd130, 8'd146, 8'd86, 8'd154, 8'd160, 8'd113, 8'd171, 8'd140, 8'd154, 8'd94, 8'd80, 8'd116, 8'd151, 8'd94, 8'd121, 8'd160, 8'd156, 8'd84, 8'd120, 8'd100, 8'd83, 8'd68, 8'd140, 8'd139, 8'd119, 8'd114, 8'd153, 8'd132, 8'd162, 8'd150, 8'd167, 8'd85, 8'd167, 8'd93, 8'd67, 8'd111, 8'd98, 8'd121, 8'd92, 8'd121, 8'd152, 8'd108, 8'd157, 8'd110, 8'd138, 8'd81, 8'd177, 8'd176, 8'd135, 8'd124, 8'd94, 8'd120, 8'd87, 8'd98, 8'd70, 8'd85, 8'd120, 8'd119, 8'd127, 8'd135, 8'd128, 8'd123, 8'd143, 8'd113, 8'd164, 8'd160, 8'd91, 8'd137, 8'd154, 8'd91, 8'd95, 8'd146, 8'd159, 8'd96, 8'd119, 8'd152, 8'd136, 8'd135, 8'd156, 8'd79, 8'd78, 8'd123, 8'd136, 8'd80, 8'd103, 8'd129, 8'd139, 8'd114, 8'd83, 8'd82, 8'd83, 8'd175, 8'd152, 8'd152, 8'd169, 8'd112, 8'd87, 8'd88, 8'd91, 8'd148, 8'd101, 8'd75, 8'd137, 8'd126, 8'd122, 8'd86, 8'd145, 8'd130, 8'd111, 8'd155, 8'd170, 8'd102, 8'd108, 8'd152, 8'd121, 8'd153, 8'd120, 8'd148, 8'd84, 8'd124, 8'd167, 8'd127, 8'd159, 8'd117, 8'd90, 8'd63, 8'd91, 8'd98, 8'd130, 8'd120, 8'd150, 8'd143, 8'd185, 8'd166, 8'd138, 8'd92, 8'd105, 8'd164, 8'd132, 8'd79, 8'd80, 8'd105, 8'd80, 8'd178, 8'd111, 8'd102, 8'd151, 8'd169, 8'd167, 8'd78, 8'd148, 8'd126, 8'd154, 8'd118, 8'd94, 8'd85, 8'd129, 8'd188, 8'd115, 8'd101, 8'd123, 8'd178, 8'd100, 8'd125, 8'd142, 8'd147, 8'd71, 8'd144, 8'd135, 8'd128, 8'd90, 8'd165, 8'd84, 8'd81, 8'd161, 8'd131, 8'd137, 8'd94, 8'd164, 8'd102, 8'd85, 8'd72, 8'd114, 8'd162, 8'd155, 8'd159, 8'd131, 8'd146, 8'd136, 8'd176, 8'd116, 8'd165, 8'd128, 8'd75, 8'd83, 8'd106, 8'd96, 8'd153, 8'd113, 8'd111, 8'd124, 8'd153, 8'd126, 8'd138, 8'd80, 8'd83, 8'd169, 8'd136, 8'd59, 8'd154, 8'd90, 8'd100, 8'd133, 8'd109, 8'd129, 8'd169, 8'd116, 8'd183, 8'd168, 8'd99, 8'd86, 8'd53, 8'd156, 8'd146, 8'd115, 8'd180, 8'd141, 8'd120, 8'd67, 8'd153, 8'd132, 8'd172, 8'd147, 8'd140, 8'd127, 8'd165, 8'd131, 8'd80, 8'd106, 8'd112, 8'd157, 8'd137, 8'd122, 8'd116, 8'd166, 8'd134, 8'd100, 8'd71, 8'd93, 8'd116, 8'd110, 8'd101, 8'd159, 8'd117, 8'd191, 8'd136, 8'd91, 8'd147, 8'd150, 8'd111, 8'd103, 8'd170, 8'd169, 8'd149, 8'd121, 8'd127, 8'd107, 8'd153, 8'd135, 8'd117, 8'd107, 8'd141, 8'd146, 8'd156, 8'd114, 8'd126, 8'd95, 8'd106, 8'd150, 8'd205, 8'd167, 8'd169, 8'd96, 8'd136, 8'd147, 8'd160, 8'd89, 8'd160, 8'd109, 8'd147, 8'd78, 8'd54, 8'd78, 8'd157, 8'd94, 8'd122, 8'd93, 8'd123, 8'd100, 8'd156, 8'd90, 8'd85, 8'd134, 8'd126, 8'd152, 8'd180, 8'd194, 8'd126, 8'd179, 8'd92, 8'd158, 8'd111, 8'd86, 8'd117, 8'd105, 8'd61, 8'd133, 8'd117, 8'd91, 8'd83, 8'd118, 8'd169, 8'd127, 8'd100, 8'd157, 8'd142, 8'd87, 8'd134, 8'd86, 8'd94, 8'd133, 8'd118, 8'd175, 8'd170, 8'd134, 8'd167, 8'd126, 8'd101, 8'd98, 8'd93, 8'd71, 8'd116, 8'd114, 8'd107, 8'd106, 8'd69, 8'd106, 8'd158, 8'd56, 8'd154, 8'd196, 8'd195, 8'd131, 8'd158, 8'd129, 8'd127, 8'd119, 8'd164, 8'd106, 8'd182, 8'd96, 8'd142, 8'd194, 8'd109, 8'd84, 8'd165, 8'd166, 8'd84, 8'd104, 8'd95, 8'd128, 8'd60, 8'd58, 8'd60, 8'd95, 8'd72, 8'd117, 8'd153, 8'd199, 8'd204, 8'd161, 8'd151, 8'd144, 8'd105, 8'd149, 8'd88, 8'd111, 8'd158, 8'd154, 8'd140, 8'd171, 8'd153, 8'd125, 8'd120, 8'd81, 8'd106, 8'd73, 8'd107, 8'd149, 8'd85, 8'd79, 8'd126, 8'd73, 8'd110, 8'd85, 8'd42, 8'd108, 8'd145, 8'd144, 8'd181, 8'd155, 8'd80, 8'd73, 8'd83, 8'd130, 8'd72, 8'd73, 8'd91, 8'd118, 8'd140, 8'd103, 8'd163, 8'd97, 8'd79, 8'd167, 8'd109, 8'd62, 8'd69, 8'd79, 8'd56, 8'd109, 8'd150, 8'd95, 8'd66, 8'd130, 8'd145, 8'd118, 8'd93, 8'd155, 8'd95, 8'd152, 8'd138, 8'd86, 8'd115, 8'd117, 8'd159, 8'd110, 8'd138, 8'd97, 8'd105, 8'd147, 8'd108, 8'd154, 8'd146, 8'd133, 8'd136, 8'd114, 8'd97, 8'd108, 8'd90, 8'd69, 8'd66, 8'd67, 8'd57, 8'd129, 8'd116, 8'd134, 8'd89, 8'd71, 8'd104, 8'd106, 8'd158, 8'd128, 8'd160, 8'd98, 8'd112, 8'd94, 8'd94, 8'd87, 8'd113, 8'd171, 8'd121, 8'd117, 8'd67, 8'd135, 8'd75, 8'd79, 8'd139, 8'd82, 8'd51, 8'd108, 8'd94, 8'd125, 8'd121, 8'd104, 8'd72, 8'd72, 8'd111, 8'd144, 8'd166, 8'd96, 8'd94, 8'd138, 8'd101, 8'd136, 8'd128, 8'd136, 8'd67, 8'd152, 8'd89, 8'd125, 8'd95, 8'd92, 8'd98, 8'd133, 8'd94, 8'd62, 8'd113, 8'd117, 8'd148, 8'd135, 8'd95, 8'd131, 8'd84, 8'd106, 8'd110, 8'd130, 8'd109, 8'd124, 8'd129, 8'd162, 8'd106, 8'd98, 8'd86, 8'd106, 8'd119, 8'd117, 8'd141, 8'd150, 8'd94, 8'd64, 8'd94, 8'd167, 8'd120, 8'd119, 8'd102, 8'd141, 8'd67, 8'd95, 8'd154, 8'd65, 8'd141, 8'd172, 8'd167, 8'd123, 8'd119, 8'd130, 8'd152, 8'd160, 8'd85, 8'd170, 8'd100, 8'd133, 8'd70, 8'd85, 8'd135, 8'd115, 8'd142, 8'd114, 8'd105, 8'd169, 8'd161, 8'd95, 8'd139, 8'd98, 8'd56, 8'd92, 8'd142, 8'd89, 8'd113, 8'd100, 8'd112, 8'd143, 8'd180, 8'd100, 8'd143, 8'd154, 8'd92, 8'd155, 8'd115, 8'd165, 8'd145, 8'd115, 8'd143, 8'd137, 8'd150, 8'd101, 8'd163, 8'd100, 8'd113, 8'd168, 8'd96, 8'd128, 8'd155, 8'd123, 8'd89, 8'd147, 8'd166, 8'd125, 8'd135, 8'd84, 8'd127, 8'd157, 8'd132, 8'd171, 8'd119, 8'd154, 8'd100, 8'd185, 8'd126, 8'd122, 8'd177, 8'd174, 8'd141, 8'd148, 8'd106, 8'd73, 8'd155, 8'd91, 8'd130, 8'd164, 8'd175, 8'd120, 8'd93, 8'd83, 8'd105, 8'd133, 8'd152, 8'd159, 8'd171, 8'd175, 8'd155, 8'd192, 8'd146, 8'd192, 8'd130, 8'd160, 8'd159, 8'd138, 8'd88, 8'd155, 8'd138, 8'd149, 8'd87, 8'd98, 8'd113, 8'd103, 8'd153, 8'd109, 8'd177, 8'd113, 8'd163, 8'd118, 8'd97, 8'd105, 8'd163, 8'd122, 8'd147, 8'd205, 8'd116, 8'd122, 8'd170, 8'd188, 8'd109, 8'd107, 8'd181, 8'd118, 8'd106, 8'd92, 8'd92, 8'd83, 8'd80, 8'd127, 8'd122, 8'd97, 8'd77, 8'd140, 8'd104, 8'd167, 8'd150, 8'd133, 8'd97, 8'd129, 8'd160, 8'd99, 8'd188, 8'd145, 8'd138, 8'd141, 8'd108, 8'd115, 8'd190, 8'd85, 8'd96, 8'd110, 8'd84, 8'd110, 8'd98, 8'd141, 8'd165, 8'd78, 8'd131, 8'd164, 8'd155, 8'd72, 8'd124, 8'd123, 8'd86, 8'd119, 8'd71, 8'd78, 8'd77, 8'd94, 8'd142, 8'd101, 8'd130, 8'd124, 8'd138, 8'd106, 8'd164, 8'd168, 8'd109, 8'd72, 8'd163, 8'd142, 8'd98, 8'd146, 8'd77, 8'd71})
) cell_0_46 (
    .clk(clk),
    .input_index(index_0_45_46),
    .input_value(value_0_45_46),
    .input_result(result_0_45_46),
    .input_enable(enable_0_45_46),
    .output_index(index_0_46_47),
    .output_value(value_0_46_47),
    .output_result(result_0_46_47),
    .output_enable(enable_0_46_47)
);

wire [10-1:0] index_0_47_48;
wire [`DATA_WIDTH-1:0] value_0_47_48;
wire [`DATA_WIDTH*4:0] result_0_47_48;
wire enable_0_47_48;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd138, 8'd78, 8'd131, 8'd98, 8'd166, 8'd90, 8'd125, 8'd102, 8'd164, 8'd145, 8'd178, 8'd174, 8'd195, 8'd180, 8'd195, 8'd88, 8'd113, 8'd183, 8'd108, 8'd93, 8'd119, 8'd100, 8'd86, 8'd89, 8'd166, 8'd146, 8'd153, 8'd109, 8'd106, 8'd161, 8'd92, 8'd127, 8'd144, 8'd171, 8'd166, 8'd152, 8'd178, 8'd143, 8'd183, 8'd171, 8'd117, 8'd125, 8'd126, 8'd114, 8'd171, 8'd142, 8'd167, 8'd142, 8'd173, 8'd82, 8'd94, 8'd100, 8'd96, 8'd163, 8'd155, 8'd99, 8'd112, 8'd145, 8'd166, 8'd120, 8'd87, 8'd111, 8'd111, 8'd75, 8'd114, 8'd140, 8'd70, 8'd133, 8'd53, 8'd141, 8'd80, 8'd152, 8'd62, 8'd48, 8'd128, 8'd119, 8'd98, 8'd100, 8'd117, 8'd108, 8'd167, 8'd105, 8'd101, 8'd112, 8'd143, 8'd180, 8'd177, 8'd149, 8'd96, 8'd90, 8'd79, 8'd101, 8'd130, 8'd141, 8'd52, 8'd70, 8'd85, 8'd100, 8'd95, 8'd143, 8'd130, 8'd53, 8'd83, 8'd83, 8'd124, 8'd162, 8'd82, 8'd77, 8'd121, 8'd158, 8'd154, 8'd85, 8'd71, 8'd87, 8'd152, 8'd156, 8'd144, 8'd140, 8'd69, 8'd82, 8'd86, 8'd85, 8'd142, 8'd126, 8'd143, 8'd91, 8'd131, 8'd125, 8'd85, 8'd136, 8'd64, 8'd87, 8'd153, 8'd129, 8'd98, 8'd72, 8'd124, 8'd155, 8'd81, 8'd136, 8'd161, 8'd160, 8'd144, 8'd93, 8'd138, 8'd95, 8'd125, 8'd102, 8'd93, 8'd122, 8'd162, 8'd136, 8'd127, 8'd156, 8'd126, 8'd124, 8'd138, 8'd129, 8'd149, 8'd164, 8'd99, 8'd92, 8'd174, 8'd88, 8'd123, 8'd61, 8'd145, 8'd100, 8'd158, 8'd172, 8'd79, 8'd155, 8'd139, 8'd51, 8'd59, 8'd106, 8'd108, 8'd163, 8'd121, 8'd69, 8'd148, 8'd132, 8'd81, 8'd93, 8'd135, 8'd180, 8'd122, 8'd137, 8'd111, 8'd83, 8'd148, 8'd61, 8'd89, 8'd90, 8'd84, 8'd111, 8'd83, 8'd160, 8'd158, 8'd91, 8'd113, 8'd122, 8'd136, 8'd118, 8'd61, 8'd145, 8'd91, 8'd63, 8'd77, 8'd89, 8'd120, 8'd127, 8'd107, 8'd126, 8'd82, 8'd124, 8'd103, 8'd64, 8'd94, 8'd74, 8'd104, 8'd83, 8'd169, 8'd103, 8'd176, 8'd160, 8'd93, 8'd151, 8'd150, 8'd108, 8'd79, 8'd142, 8'd98, 8'd146, 8'd121, 8'd124, 8'd103, 8'd159, 8'd179, 8'd171, 8'd166, 8'd131, 8'd154, 8'd90, 8'd131, 8'd77, 8'd72, 8'd121, 8'd57, 8'd124, 8'd173, 8'd93, 8'd163, 8'd145, 8'd148, 8'd116, 8'd106, 8'd147, 8'd101, 8'd147, 8'd60, 8'd102, 8'd85, 8'd149, 8'd80, 8'd91, 8'd139, 8'd194, 8'd140, 8'd142, 8'd127, 8'd109, 8'd128, 8'd129, 8'd79, 8'd139, 8'd57, 8'd127, 8'd133, 8'd180, 8'd89, 8'd116, 8'd163, 8'd111, 8'd118, 8'd115, 8'd96, 8'd108, 8'd65, 8'd123, 8'd112, 8'd153, 8'd121, 8'd138, 8'd181, 8'd102, 8'd160, 8'd141, 8'd173, 8'd124, 8'd131, 8'd68, 8'd118, 8'd123, 8'd56, 8'd124, 8'd162, 8'd153, 8'd175, 8'd152, 8'd97, 8'd146, 8'd164, 8'd107, 8'd90, 8'd141, 8'd119, 8'd132, 8'd126, 8'd72, 8'd137, 8'd148, 8'd174, 8'd161, 8'd115, 8'd132, 8'd136, 8'd156, 8'd101, 8'd145, 8'd119, 8'd106, 8'd114, 8'd158, 8'd143, 8'd160, 8'd119, 8'd85, 8'd112, 8'd120, 8'd162, 8'd112, 8'd154, 8'd131, 8'd100, 8'd85, 8'd138, 8'd145, 8'd116, 8'd110, 8'd130, 8'd52, 8'd110, 8'd115, 8'd125, 8'd170, 8'd110, 8'd105, 8'd156, 8'd82, 8'd88, 8'd172, 8'd89, 8'd153, 8'd112, 8'd102, 8'd121, 8'd132, 8'd155, 8'd115, 8'd150, 8'd79, 8'd92, 8'd104, 8'd133, 8'd68, 8'd80, 8'd70, 8'd115, 8'd66, 8'd110, 8'd48, 8'd93, 8'd116, 8'd105, 8'd121, 8'd78, 8'd122, 8'd110, 8'd152, 8'd104, 8'd65, 8'd125, 8'd90, 8'd99, 8'd149, 8'd118, 8'd149, 8'd120, 8'd90, 8'd121, 8'd60, 8'd55, 8'd144, 8'd158, 8'd80, 8'd85, 8'd111, 8'd104, 8'd132, 8'd125, 8'd71, 8'd147, 8'd93, 8'd157, 8'd148, 8'd141, 8'd181, 8'd108, 8'd95, 8'd172, 8'd109, 8'd135, 8'd119, 8'd139, 8'd132, 8'd166, 8'd146, 8'd159, 8'd105, 8'd89, 8'd122, 8'd85, 8'd67, 8'd96, 8'd90, 8'd104, 8'd131, 8'd77, 8'd77, 8'd106, 8'd142, 8'd113, 8'd117, 8'd146, 8'd99, 8'd163, 8'd97, 8'd129, 8'd105, 8'd26, 8'd95, 8'd132, 8'd171, 8'd155, 8'd147, 8'd89, 8'd164, 8'd164, 8'd154, 8'd146, 8'd165, 8'd84, 8'd136, 8'd151, 8'd148, 8'd74, 8'd151, 8'd160, 8'd140, 8'd92, 8'd159, 8'd128, 8'd119, 8'd156, 8'd169, 8'd104, 8'd56, 8'd59, 8'd116, 8'd80, 8'd89, 8'd113, 8'd157, 8'd128, 8'd115, 8'd95, 8'd170, 8'd134, 8'd99, 8'd85, 8'd134, 8'd166, 8'd136, 8'd129, 8'd66, 8'd116, 8'd163, 8'd140, 8'd117, 8'd179, 8'd172, 8'd95, 8'd93, 8'd73, 8'd126, 8'd63, 8'd127, 8'd86, 8'd81, 8'd149, 8'd94, 8'd146, 8'd81, 8'd143, 8'd194, 8'd103, 8'd91, 8'd84, 8'd116, 8'd146, 8'd154, 8'd86, 8'd136, 8'd79, 8'd110, 8'd155, 8'd131, 8'd123, 8'd160, 8'd135, 8'd139, 8'd106, 8'd72, 8'd85, 8'd121, 8'd94, 8'd149, 8'd107, 8'd96, 8'd112, 8'd135, 8'd99, 8'd98, 8'd155, 8'd107, 8'd147, 8'd157, 8'd125, 8'd95, 8'd158, 8'd84, 8'd159, 8'd92, 8'd165, 8'd146, 8'd167, 8'd132, 8'd157, 8'd168, 8'd148, 8'd59, 8'd65, 8'd75, 8'd131, 8'd129, 8'd136, 8'd132, 8'd90, 8'd93, 8'd68, 8'd122, 8'd104, 8'd115, 8'd145, 8'd95, 8'd101, 8'd103, 8'd91, 8'd89, 8'd97, 8'd154, 8'd135, 8'd161, 8'd166, 8'd184, 8'd111, 8'd112, 8'd84, 8'd119, 8'd63, 8'd85, 8'd125, 8'd159, 8'd97, 8'd75, 8'd74, 8'd91, 8'd96, 8'd125, 8'd90, 8'd136, 8'd151, 8'd110, 8'd128, 8'd142, 8'd87, 8'd134, 8'd115, 8'd109, 8'd123, 8'd93, 8'd142, 8'd85, 8'd153, 8'd106, 8'd164, 8'd112, 8'd106, 8'd133, 8'd76, 8'd153, 8'd136, 8'd173, 8'd144, 8'd77, 8'd129, 8'd105, 8'd129, 8'd93, 8'd99, 8'd71, 8'd77, 8'd100, 8'd118, 8'd105, 8'd81, 8'd102, 8'd86, 8'd155, 8'd159, 8'd99, 8'd113, 8'd159, 8'd134, 8'd118, 8'd143, 8'd110, 8'd123, 8'd95, 8'd148, 8'd100, 8'd148, 8'd140, 8'd146, 8'd109, 8'd95, 8'd98, 8'd131, 8'd120, 8'd131, 8'd147, 8'd68, 8'd149, 8'd161, 8'd97, 8'd165, 8'd155, 8'd69, 8'd93, 8'd86, 8'd74, 8'd95, 8'd75, 8'd167, 8'd171, 8'd92, 8'd85, 8'd149, 8'd97, 8'd106, 8'd101, 8'd80, 8'd90, 8'd116, 8'd148, 8'd102, 8'd123, 8'd115, 8'd150, 8'd164, 8'd170, 8'd109, 8'd106, 8'd100, 8'd164, 8'd98, 8'd103, 8'd73, 8'd95, 8'd140, 8'd116, 8'd173, 8'd119, 8'd129, 8'd92, 8'd123, 8'd174, 8'd137, 8'd160, 8'd130, 8'd181, 8'd148, 8'd197, 8'd126, 8'd137, 8'd156, 8'd163, 8'd195, 8'd158, 8'd171, 8'd163, 8'd81, 8'd168, 8'd87, 8'd121, 8'd168, 8'd94, 8'd88, 8'd108, 8'd128, 8'd151, 8'd94, 8'd171, 8'd129, 8'd128, 8'd123, 8'd182, 8'd173, 8'd186, 8'd125, 8'd136, 8'd147, 8'd167, 8'd104, 8'd122, 8'd108, 8'd95, 8'd127, 8'd183, 8'd175, 8'd143, 8'd135, 8'd163, 8'd86, 8'd159, 8'd94, 8'd112, 8'd77, 8'd111, 8'd137, 8'd87, 8'd130, 8'd98, 8'd133, 8'd152, 8'd88, 8'd122, 8'd102, 8'd118, 8'd111, 8'd118, 8'd102, 8'd80, 8'd111, 8'd105, 8'd142, 8'd104, 8'd110, 8'd154, 8'd128, 8'd115, 8'd110, 8'd91})
) cell_0_47 (
    .clk(clk),
    .input_index(index_0_46_47),
    .input_value(value_0_46_47),
    .input_result(result_0_46_47),
    .input_enable(enable_0_46_47),
    .output_index(index_0_47_48),
    .output_value(value_0_47_48),
    .output_result(result_0_47_48),
    .output_enable(enable_0_47_48)
);

wire [10-1:0] index_0_48_49;
wire [`DATA_WIDTH-1:0] value_0_48_49;
wire [`DATA_WIDTH*4:0] result_0_48_49;
wire enable_0_48_49;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd81, 8'd148, 8'd81, 8'd130, 8'd112, 8'd75, 8'd100, 8'd80, 8'd73, 8'd98, 8'd126, 8'd130, 8'd145, 8'd119, 8'd94, 8'd113, 8'd89, 8'd107, 8'd151, 8'd93, 8'd132, 8'd89, 8'd123, 8'd81, 8'd82, 8'd93, 8'd143, 8'd86, 8'd92, 8'd138, 8'd94, 8'd152, 8'd104, 8'd100, 8'd69, 8'd108, 8'd136, 8'd72, 8'd106, 8'd110, 8'd66, 8'd100, 8'd105, 8'd129, 8'd137, 8'd93, 8'd113, 8'd107, 8'd158, 8'd157, 8'd145, 8'd164, 8'd153, 8'd87, 8'd106, 8'd152, 8'd128, 8'd116, 8'd113, 8'd112, 8'd96, 8'd114, 8'd144, 8'd142, 8'd173, 8'd151, 8'd65, 8'd111, 8'd97, 8'd150, 8'd108, 8'd152, 8'd96, 8'd160, 8'd135, 8'd126, 8'd147, 8'd112, 8'd143, 8'd60, 8'd150, 8'd125, 8'd116, 8'd80, 8'd79, 8'd67, 8'd119, 8'd121, 8'd149, 8'd157, 8'd151, 8'd192, 8'd160, 8'd170, 8'd170, 8'd81, 8'd82, 8'd108, 8'd73, 8'd119, 8'd145, 8'd144, 8'd141, 8'd143, 8'd168, 8'd77, 8'd146, 8'd58, 8'd91, 8'd107, 8'd132, 8'd128, 8'd74, 8'd110, 8'd100, 8'd168, 8'd112, 8'd142, 8'd113, 8'd160, 8'd173, 8'd85, 8'd147, 8'd168, 8'd148, 8'd125, 8'd138, 8'd156, 8'd133, 8'd143, 8'd147, 8'd138, 8'd87, 8'd81, 8'd147, 8'd48, 8'd144, 8'd146, 8'd129, 8'd147, 8'd161, 8'd160, 8'd68, 8'd147, 8'd122, 8'd135, 8'd154, 8'd100, 8'd106, 8'd151, 8'd99, 8'd123, 8'd75, 8'd83, 8'd111, 8'd70, 8'd125, 8'd150, 8'd98, 8'd70, 8'd115, 8'd135, 8'd134, 8'd81, 8'd72, 8'd129, 8'd156, 8'd145, 8'd99, 8'd139, 8'd70, 8'd166, 8'd162, 8'd146, 8'd112, 8'd157, 8'd93, 8'd119, 8'd156, 8'd90, 8'd119, 8'd106, 8'd138, 8'd125, 8'd71, 8'd128, 8'd62, 8'd106, 8'd98, 8'd61, 8'd147, 8'd143, 8'd42, 8'd146, 8'd152, 8'd113, 8'd95, 8'd132, 8'd62, 8'd101, 8'd144, 8'd60, 8'd60, 8'd122, 8'd87, 8'd146, 8'd80, 8'd73, 8'd115, 8'd121, 8'd38, 8'd124, 8'd105, 8'd19, 8'd30, 8'd76, 8'd69, 8'd71, 8'd59, 8'd52, 8'd53, 8'd99, 8'd81, 8'd158, 8'd76, 8'd127, 8'd124, 8'd74, 8'd103, 8'd80, 8'd111, 8'd115, 8'd107, 8'd77, 8'd96, 8'd117, 8'd126, 8'd99, 8'd141, 8'd72, 8'd55, 8'd91, 8'd125, 8'd55, 8'd149, 8'd149, 8'd70, 8'd54, 8'd56, 8'd65, 8'd126, 8'd82, 8'd117, 8'd136, 8'd115, 8'd88, 8'd102, 8'd115, 8'd96, 8'd148, 8'd87, 8'd142, 8'd122, 8'd75, 8'd167, 8'd110, 8'd91, 8'd136, 8'd127, 8'd122, 8'd78, 8'd140, 8'd105, 8'd62, 8'd91, 8'd107, 8'd98, 8'd119, 8'd67, 8'd152, 8'd127, 8'd102, 8'd30, 8'd29, 8'd52, 8'd58, 8'd72, 8'd146, 8'd89, 8'd68, 8'd98, 8'd116, 8'd125, 8'd143, 8'd150, 8'd89, 8'd110, 8'd154, 8'd142, 8'd186, 8'd90, 8'd104, 8'd72, 8'd44, 8'd81, 8'd123, 8'd80, 8'd164, 8'd92, 8'd106, 8'd64, 8'd80, 8'd60, 8'd132, 8'd111, 8'd123, 8'd100, 8'd90, 8'd96, 8'd113, 8'd97, 8'd164, 8'd90, 8'd112, 8'd115, 8'd131, 8'd88, 8'd170, 8'd129, 8'd89, 8'd137, 8'd130, 8'd56, 8'd104, 8'd134, 8'd141, 8'd66, 8'd156, 8'd128, 8'd108, 8'd63, 8'd54, 8'd95, 8'd101, 8'd145, 8'd166, 8'd165, 8'd139, 8'd123, 8'd72, 8'd126, 8'd101, 8'd168, 8'd98, 8'd137, 8'd129, 8'd158, 8'd140, 8'd138, 8'd118, 8'd163, 8'd70, 8'd73, 8'd111, 8'd68, 8'd93, 8'd127, 8'd116, 8'd63, 8'd152, 8'd93, 8'd91, 8'd118, 8'd144, 8'd119, 8'd194, 8'd94, 8'd148, 8'd169, 8'd121, 8'd96, 8'd174, 8'd178, 8'd126, 8'd164, 8'd117, 8'd168, 8'd111, 8'd90, 8'd112, 8'd125, 8'd120, 8'd121, 8'd99, 8'd70, 8'd118, 8'd98, 8'd139, 8'd140, 8'd124, 8'd106, 8'd151, 8'd153, 8'd191, 8'd116, 8'd184, 8'd91, 8'd144, 8'd165, 8'd162, 8'd180, 8'd121, 8'd106, 8'd109, 8'd137, 8'd92, 8'd135, 8'd88, 8'd87, 8'd89, 8'd140, 8'd66, 8'd55, 8'd103, 8'd130, 8'd116, 8'd114, 8'd120, 8'd96, 8'd121, 8'd104, 8'd179, 8'd190, 8'd119, 8'd131, 8'd138, 8'd141, 8'd170, 8'd158, 8'd166, 8'd152, 8'd185, 8'd165, 8'd140, 8'd150, 8'd108, 8'd102, 8'd154, 8'd110, 8'd105, 8'd64, 8'd34, 8'd90, 8'd115, 8'd109, 8'd120, 8'd165, 8'd158, 8'd110, 8'd184, 8'd153, 8'd62, 8'd74, 8'd166, 8'd148, 8'd171, 8'd175, 8'd160, 8'd175, 8'd116, 8'd137, 8'd81, 8'd107, 8'd60, 8'd127, 8'd66, 8'd92, 8'd30, 8'd106, 8'd81, 8'd110, 8'd134, 8'd131, 8'd135, 8'd153, 8'd83, 8'd120, 8'd71, 8'd65, 8'd43, 8'd103, 8'd118, 8'd138, 8'd160, 8'd100, 8'd103, 8'd105, 8'd103, 8'd120, 8'd126, 8'd65, 8'd130, 8'd66, 8'd95, 8'd81, 8'd131, 8'd122, 8'd79, 8'd121, 8'd155, 8'd118, 8'd94, 8'd103, 8'd166, 8'd128, 8'd81, 8'd129, 8'd55, 8'd115, 8'd106, 8'd68, 8'd94, 8'd153, 8'd78, 8'd98, 8'd133, 8'd61, 8'd73, 8'd81, 8'd64, 8'd70, 8'd71, 8'd82, 8'd75, 8'd118, 8'd100, 8'd115, 8'd94, 8'd107, 8'd101, 8'd84, 8'd168, 8'd120, 8'd92, 8'd103, 8'd110, 8'd114, 8'd69, 8'd58, 8'd145, 8'd141, 8'd71, 8'd140, 8'd100, 8'd50, 8'd90, 8'd79, 8'd75, 8'd64, 8'd138, 8'd77, 8'd111, 8'd131, 8'd94, 8'd141, 8'd143, 8'd90, 8'd130, 8'd171, 8'd146, 8'd164, 8'd82, 8'd89, 8'd147, 8'd116, 8'd113, 8'd118, 8'd77, 8'd125, 8'd61, 8'd79, 8'd127, 8'd115, 8'd52, 8'd79, 8'd143, 8'd123, 8'd131, 8'd65, 8'd85, 8'd142, 8'd160, 8'd112, 8'd105, 8'd111, 8'd122, 8'd126, 8'd102, 8'd91, 8'd109, 8'd145, 8'd121, 8'd105, 8'd90, 8'd115, 8'd112, 8'd88, 8'd93, 8'd113, 8'd100, 8'd125, 8'd141, 8'd104, 8'd132, 8'd118, 8'd76, 8'd124, 8'd120, 8'd76, 8'd150, 8'd88, 8'd126, 8'd61, 8'd134, 8'd100, 8'd105, 8'd70, 8'd107, 8'd110, 8'd144, 8'd67, 8'd97, 8'd78, 8'd74, 8'd123, 8'd117, 8'd70, 8'd120, 8'd97, 8'd160, 8'd71, 8'd105, 8'd105, 8'd132, 8'd157, 8'd133, 8'd110, 8'd106, 8'd162, 8'd148, 8'd99, 8'd106, 8'd125, 8'd117, 8'd118, 8'd85, 8'd123, 8'd87, 8'd86, 8'd123, 8'd28, 8'd124, 8'd112, 8'd70, 8'd145, 8'd120, 8'd83, 8'd154, 8'd120, 8'd130, 8'd136, 8'd146, 8'd115, 8'd79, 8'd136, 8'd48, 8'd75, 8'd96, 8'd95, 8'd102, 8'd43, 8'd103, 8'd68, 8'd53, 8'd7, 8'd18, 8'd0, 8'd52, 8'd33, 8'd40, 8'd112, 8'd92, 8'd56, 8'd144, 8'd66, 8'd70, 8'd127, 8'd108, 8'd82, 8'd168, 8'd120, 8'd140, 8'd82, 8'd144, 8'd135, 8'd67, 8'd116, 8'd67, 8'd42, 8'd43, 8'd52, 8'd101, 8'd101, 8'd106, 8'd35, 8'd48, 8'd105, 8'd48, 8'd64, 8'd75, 8'd68, 8'd133, 8'd119, 8'd81, 8'd108, 8'd118, 8'd161, 8'd142, 8'd107, 8'd95, 8'd95, 8'd115, 8'd76, 8'd70, 8'd82, 8'd124, 8'd75, 8'd60, 8'd118, 8'd102, 8'd142, 8'd143, 8'd73, 8'd131, 8'd132, 8'd98, 8'd52, 8'd84, 8'd84, 8'd82, 8'd75, 8'd107, 8'd154, 8'd130, 8'd127, 8'd122, 8'd153, 8'd126, 8'd75, 8'd76, 8'd148, 8'd99, 8'd110, 8'd129, 8'd137, 8'd135, 8'd116, 8'd131, 8'd90, 8'd159, 8'd72, 8'd91, 8'd156, 8'd149, 8'd141, 8'd162, 8'd151, 8'd147, 8'd111, 8'd160, 8'd128, 8'd158, 8'd127, 8'd155})
) cell_0_48 (
    .clk(clk),
    .input_index(index_0_47_48),
    .input_value(value_0_47_48),
    .input_result(result_0_47_48),
    .input_enable(enable_0_47_48),
    .output_index(index_0_48_49),
    .output_value(value_0_48_49),
    .output_result(result_0_48_49),
    .output_enable(enable_0_48_49)
);

wire [10-1:0] index_0_49_50;
wire [`DATA_WIDTH-1:0] value_0_49_50;
wire [`DATA_WIDTH*4:0] result_0_49_50;
wire enable_0_49_50;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd154, 8'd120, 8'd76, 8'd138, 8'd59, 8'd155, 8'd152, 8'd160, 8'd74, 8'd104, 8'd86, 8'd77, 8'd129, 8'd143, 8'd136, 8'd80, 8'd104, 8'd136, 8'd130, 8'd131, 8'd165, 8'd104, 8'd87, 8'd93, 8'd162, 8'd162, 8'd98, 8'd86, 8'd130, 8'd85, 8'd100, 8'd124, 8'd154, 8'd140, 8'd167, 8'd155, 8'd82, 8'd132, 8'd164, 8'd91, 8'd115, 8'd108, 8'd123, 8'd119, 8'd106, 8'd139, 8'd121, 8'd90, 8'd91, 8'd158, 8'd124, 8'd139, 8'd138, 8'd110, 8'd151, 8'd114, 8'd134, 8'd91, 8'd109, 8'd77, 8'd90, 8'd107, 8'd118, 8'd113, 8'd105, 8'd178, 8'd121, 8'd105, 8'd151, 8'd109, 8'd146, 8'd79, 8'd145, 8'd123, 8'd162, 8'd159, 8'd144, 8'd77, 8'd76, 8'd148, 8'd68, 8'd117, 8'd77, 8'd91, 8'd118, 8'd142, 8'd101, 8'd101, 8'd116, 8'd187, 8'd134, 8'd158, 8'd124, 8'd137, 8'd109, 8'd106, 8'd167, 8'd162, 8'd91, 8'd73, 8'd115, 8'd90, 8'd138, 8'd106, 8'd98, 8'd143, 8'd104, 8'd61, 8'd78, 8'd87, 8'd97, 8'd115, 8'd70, 8'd144, 8'd74, 8'd128, 8'd171, 8'd101, 8'd134, 8'd124, 8'd134, 8'd96, 8'd124, 8'd105, 8'd103, 8'd141, 8'd103, 8'd156, 8'd135, 8'd85, 8'd149, 8'd74, 8'd78, 8'd94, 8'd112, 8'd90, 8'd125, 8'd153, 8'd86, 8'd71, 8'd165, 8'd69, 8'd138, 8'd96, 8'd113, 8'd115, 8'd115, 8'd111, 8'd72, 8'd78, 8'd87, 8'd152, 8'd127, 8'd116, 8'd150, 8'd169, 8'd72, 8'd70, 8'd99, 8'd80, 8'd154, 8'd127, 8'd82, 8'd73, 8'd153, 8'd125, 8'd127, 8'd121, 8'd93, 8'd133, 8'd153, 8'd97, 8'd145, 8'd197, 8'd179, 8'd86, 8'd103, 8'd164, 8'd116, 8'd82, 8'd106, 8'd162, 8'd145, 8'd143, 8'd97, 8'd98, 8'd141, 8'd119, 8'd159, 8'd108, 8'd118, 8'd91, 8'd133, 8'd64, 8'd108, 8'd69, 8'd142, 8'd125, 8'd177, 8'd174, 8'd120, 8'd103, 8'd133, 8'd160, 8'd127, 8'd138, 8'd120, 8'd150, 8'd63, 8'd109, 8'd103, 8'd64, 8'd94, 8'd113, 8'd120, 8'd115, 8'd92, 8'd160, 8'd76, 8'd110, 8'd55, 8'd125, 8'd84, 8'd104, 8'd93, 8'd77, 8'd73, 8'd181, 8'd145, 8'd168, 8'd121, 8'd137, 8'd94, 8'd93, 8'd120, 8'd69, 8'd130, 8'd129, 8'd161, 8'd147, 8'd139, 8'd101, 8'd156, 8'd129, 8'd137, 8'd83, 8'd93, 8'd127, 8'd58, 8'd97, 8'd150, 8'd86, 8'd101, 8'd98, 8'd67, 8'd173, 8'd89, 8'd122, 8'd130, 8'd133, 8'd150, 8'd148, 8'd129, 8'd116, 8'd122, 8'd104, 8'd151, 8'd131, 8'd152, 8'd102, 8'd118, 8'd87, 8'd166, 8'd175, 8'd126, 8'd126, 8'd95, 8'd93, 8'd91, 8'd107, 8'd116, 8'd150, 8'd58, 8'd134, 8'd137, 8'd144, 8'd128, 8'd150, 8'd152, 8'd85, 8'd81, 8'd111, 8'd153, 8'd128, 8'd77, 8'd115, 8'd94, 8'd123, 8'd91, 8'd169, 8'd85, 8'd138, 8'd156, 8'd87, 8'd76, 8'd58, 8'd155, 8'd106, 8'd97, 8'd68, 8'd145, 8'd75, 8'd107, 8'd98, 8'd50, 8'd66, 8'd60, 8'd84, 8'd157, 8'd107, 8'd115, 8'd79, 8'd154, 8'd176, 8'd156, 8'd168, 8'd127, 8'd82, 8'd136, 8'd61, 8'd72, 8'd61, 8'd111, 8'd57, 8'd113, 8'd102, 8'd105, 8'd74, 8'd124, 8'd112, 8'd70, 8'd45, 8'd135, 8'd79, 8'd134, 8'd138, 8'd111, 8'd90, 8'd98, 8'd127, 8'd116, 8'd149, 8'd111, 8'd99, 8'd104, 8'd105, 8'd125, 8'd98, 8'd125, 8'd133, 8'd111, 8'd122, 8'd78, 8'd94, 8'd160, 8'd160, 8'd115, 8'd39, 8'd118, 8'd88, 8'd83, 8'd87, 8'd123, 8'd132, 8'd125, 8'd118, 8'd79, 8'd120, 8'd128, 8'd124, 8'd167, 8'd161, 8'd84, 8'd126, 8'd154, 8'd89, 8'd158, 8'd81, 8'd91, 8'd55, 8'd63, 8'd90, 8'd139, 8'd95, 8'd91, 8'd25, 8'd121, 8'd139, 8'd86, 8'd94, 8'd169, 8'd143, 8'd131, 8'd108, 8'd143, 8'd173, 8'd171, 8'd147, 8'd184, 8'd126, 8'd133, 8'd160, 8'd127, 8'd171, 8'd152, 8'd154, 8'd91, 8'd129, 8'd100, 8'd105, 8'd131, 8'd119, 8'd66, 8'd54, 8'd75, 8'd123, 8'd99, 8'd165, 8'd144, 8'd93, 8'd142, 8'd95, 8'd140, 8'd173, 8'd155, 8'd142, 8'd180, 8'd88, 8'd164, 8'd106, 8'd82, 8'd181, 8'd154, 8'd145, 8'd108, 8'd82, 8'd132, 8'd74, 8'd143, 8'd147, 8'd121, 8'd113, 8'd102, 8'd79, 8'd76, 8'd112, 8'd123, 8'd122, 8'd102, 8'd121, 8'd156, 8'd97, 8'd130, 8'd109, 8'd175, 8'd86, 8'd173, 8'd97, 8'd133, 8'd137, 8'd97, 8'd95, 8'd64, 8'd58, 8'd101, 8'd84, 8'd158, 8'd199, 8'd186, 8'd197, 8'd171, 8'd100, 8'd147, 8'd136, 8'd148, 8'd108, 8'd113, 8'd50, 8'd47, 8'd72, 8'd96, 8'd122, 8'd144, 8'd151, 8'd125, 8'd124, 8'd154, 8'd81, 8'd100, 8'd141, 8'd77, 8'd132, 8'd93, 8'd101, 8'd81, 8'd184, 8'd179, 8'd200, 8'd121, 8'd72, 8'd130, 8'd112, 8'd94, 8'd73, 8'd102, 8'd144, 8'd136, 8'd80, 8'd154, 8'd100, 8'd94, 8'd102, 8'd166, 8'd126, 8'd75, 8'd149, 8'd122, 8'd91, 8'd125, 8'd81, 8'd111, 8'd107, 8'd169, 8'd197, 8'd158, 8'd136, 8'd133, 8'd119, 8'd100, 8'd141, 8'd113, 8'd81, 8'd121, 8'd89, 8'd136, 8'd151, 8'd125, 8'd98, 8'd84, 8'd164, 8'd110, 8'd131, 8'd70, 8'd103, 8'd119, 8'd130, 8'd89, 8'd86, 8'd58, 8'd100, 8'd107, 8'd167, 8'd180, 8'd163, 8'd105, 8'd108, 8'd113, 8'd119, 8'd134, 8'd152, 8'd79, 8'd140, 8'd181, 8'd183, 8'd101, 8'd135, 8'd155, 8'd158, 8'd108, 8'd123, 8'd70, 8'd134, 8'd123, 8'd74, 8'd70, 8'd125, 8'd134, 8'd132, 8'd118, 8'd183, 8'd173, 8'd115, 8'd157, 8'd124, 8'd79, 8'd168, 8'd158, 8'd147, 8'd118, 8'd154, 8'd143, 8'd173, 8'd138, 8'd79, 8'd116, 8'd131, 8'd100, 8'd149, 8'd64, 8'd90, 8'd66, 8'd94, 8'd132, 8'd79, 8'd87, 8'd121, 8'd114, 8'd124, 8'd108, 8'd122, 8'd154, 8'd123, 8'd112, 8'd123, 8'd90, 8'd140, 8'd93, 8'd103, 8'd125, 8'd127, 8'd122, 8'd83, 8'd112, 8'd80, 8'd60, 8'd107, 8'd92, 8'd127, 8'd109, 8'd87, 8'd128, 8'd125, 8'd108, 8'd168, 8'd115, 8'd161, 8'd120, 8'd102, 8'd97, 8'd116, 8'd65, 8'd94, 8'd92, 8'd140, 8'd143, 8'd108, 8'd142, 8'd144, 8'd77, 8'd149, 8'd144, 8'd99, 8'd114, 8'd149, 8'd83, 8'd91, 8'd86, 8'd137, 8'd123, 8'd150, 8'd85, 8'd158, 8'd156, 8'd79, 8'd103, 8'd129, 8'd159, 8'd111, 8'd85, 8'd98, 8'd125, 8'd137, 8'd142, 8'd136, 8'd84, 8'd73, 8'd88, 8'd113, 8'd62, 8'd65, 8'd61, 8'd85, 8'd63, 8'd90, 8'd151, 8'd94, 8'd120, 8'd117, 8'd87, 8'd151, 8'd158, 8'd167, 8'd127, 8'd58, 8'd80, 8'd149, 8'd72, 8'd110, 8'd131, 8'd87, 8'd147, 8'd108, 8'd112, 8'd104, 8'd84, 8'd73, 8'd54, 8'd93, 8'd129, 8'd111, 8'd102, 8'd130, 8'd62, 8'd160, 8'd87, 8'd110, 8'd83, 8'd168, 8'd128, 8'd121, 8'd93, 8'd146, 8'd138, 8'd109, 8'd146, 8'd144, 8'd66, 8'd80, 8'd121, 8'd102, 8'd97, 8'd134, 8'd68, 8'd148, 8'd98, 8'd110, 8'd105, 8'd121, 8'd70, 8'd131, 8'd160, 8'd121, 8'd163, 8'd133, 8'd100, 8'd101, 8'd159, 8'd77, 8'd154, 8'd110, 8'd91, 8'd129, 8'd100, 8'd165, 8'd137, 8'd87, 8'd85, 8'd119, 8'd146, 8'd113, 8'd94, 8'd149, 8'd91, 8'd153, 8'd135, 8'd96, 8'd73, 8'd113, 8'd78, 8'd168, 8'd86, 8'd73, 8'd167, 8'd169})
) cell_0_49 (
    .clk(clk),
    .input_index(index_0_48_49),
    .input_value(value_0_48_49),
    .input_result(result_0_48_49),
    .input_enable(enable_0_48_49),
    .output_index(index_0_49_50),
    .output_value(value_0_49_50),
    .output_result(result_0_49_50),
    .output_enable(enable_0_49_50)
);

wire [10-1:0] index_0_50_51;
wire [`DATA_WIDTH-1:0] value_0_50_51;
wire [`DATA_WIDTH*4:0] result_0_50_51;
wire enable_0_50_51;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd72, 8'd82, 8'd119, 8'd113, 8'd70, 8'd162, 8'd84, 8'd88, 8'd162, 8'd141, 8'd168, 8'd133, 8'd150, 8'd127, 8'd136, 8'd168, 8'd119, 8'd168, 8'd110, 8'd136, 8'd171, 8'd119, 8'd134, 8'd116, 8'd84, 8'd161, 8'd86, 8'd144, 8'd110, 8'd150, 8'd110, 8'd173, 8'd85, 8'd161, 8'd184, 8'd172, 8'd200, 8'd129, 8'd201, 8'd128, 8'd185, 8'd205, 8'd196, 8'd161, 8'd177, 8'd151, 8'd110, 8'd96, 8'd182, 8'd111, 8'd98, 8'd80, 8'd131, 8'd120, 8'd140, 8'd74, 8'd162, 8'd161, 8'd110, 8'd180, 8'd78, 8'd151, 8'd168, 8'd105, 8'd169, 8'd98, 8'd139, 8'd177, 8'd115, 8'd155, 8'd176, 8'd114, 8'd120, 8'd113, 8'd170, 8'd168, 8'd117, 8'd92, 8'd118, 8'd105, 8'd72, 8'd159, 8'd129, 8'd149, 8'd80, 8'd114, 8'd143, 8'd145, 8'd126, 8'd157, 8'd134, 8'd136, 8'd101, 8'd134, 8'd148, 8'd126, 8'd146, 8'd157, 8'd157, 8'd116, 8'd86, 8'd106, 8'd120, 8'd84, 8'd125, 8'd132, 8'd60, 8'd127, 8'd149, 8'd156, 8'd162, 8'd166, 8'd91, 8'd107, 8'd161, 8'd154, 8'd189, 8'd146, 8'd116, 8'd164, 8'd140, 8'd128, 8'd66, 8'd95, 8'd112, 8'd106, 8'd138, 8'd142, 8'd123, 8'd148, 8'd149, 8'd167, 8'd184, 8'd136, 8'd177, 8'd140, 8'd172, 8'd120, 8'd163, 8'd160, 8'd165, 8'd160, 8'd173, 8'd178, 8'd199, 8'd189, 8'd169, 8'd105, 8'd178, 8'd96, 8'd167, 8'd88, 8'd97, 8'd128, 8'd76, 8'd106, 8'd180, 8'd132, 8'd202, 8'd187, 8'd125, 8'd156, 8'd192, 8'd126, 8'd142, 8'd179, 8'd76, 8'd103, 8'd132, 8'd122, 8'd170, 8'd134, 8'd183, 8'd188, 8'd110, 8'd115, 8'd135, 8'd166, 8'd155, 8'd76, 8'd66, 8'd60, 8'd72, 8'd72, 8'd165, 8'd131, 8'd145, 8'd114, 8'd180, 8'd192, 8'd132, 8'd117, 8'd142, 8'd131, 8'd165, 8'd105, 8'd113, 8'd106, 8'd130, 8'd140, 8'd135, 8'd187, 8'd151, 8'd94, 8'd137, 8'd117, 8'd156, 8'd123, 8'd96, 8'd85, 8'd109, 8'd129, 8'd158, 8'd175, 8'd124, 8'd155, 8'd179, 8'd141, 8'd170, 8'd182, 8'd156, 8'd89, 8'd124, 8'd105, 8'd131, 8'd104, 8'd196, 8'd195, 8'd199, 8'd167, 8'd133, 8'd103, 8'd116, 8'd130, 8'd157, 8'd146, 8'd80, 8'd112, 8'd102, 8'd96, 8'd117, 8'd182, 8'd158, 8'd164, 8'd173, 8'd176, 8'd115, 8'd180, 8'd105, 8'd167, 8'd111, 8'd122, 8'd139, 8'd148, 8'd122, 8'd190, 8'd124, 8'd141, 8'd127, 8'd93, 8'd92, 8'd107, 8'd110, 8'd125, 8'd79, 8'd154, 8'd95, 8'd84, 8'd124, 8'd106, 8'd134, 8'd79, 8'd81, 8'd113, 8'd140, 8'd213, 8'd210, 8'd113, 8'd117, 8'd161, 8'd113, 8'd181, 8'd176, 8'd196, 8'd141, 8'd138, 8'd89, 8'd77, 8'd64, 8'd66, 8'd109, 8'd128, 8'd67, 8'd135, 8'd75, 8'd144, 8'd58, 8'd118, 8'd124, 8'd109, 8'd125, 8'd134, 8'd198, 8'd152, 8'd144, 8'd106, 8'd100, 8'd109, 8'd114, 8'd110, 8'd208, 8'd158, 8'd116, 8'd154, 8'd161, 8'd58, 8'd128, 8'd112, 8'd64, 8'd65, 8'd75, 8'd116, 8'd125, 8'd134, 8'd91, 8'd110, 8'd35, 8'd89, 8'd62, 8'd68, 8'd91, 8'd201, 8'd190, 8'd125, 8'd126, 8'd93, 8'd133, 8'd159, 8'd149, 8'd186, 8'd55, 8'd70, 8'd54, 8'd120, 8'd141, 8'd106, 8'd125, 8'd107, 8'd124, 8'd102, 8'd142, 8'd121, 8'd32, 8'd112, 8'd42, 8'd59, 8'd118, 8'd125, 8'd141, 8'd147, 8'd125, 8'd108, 8'd98, 8'd169, 8'd168, 8'd112, 8'd127, 8'd150, 8'd106, 8'd108, 8'd102, 8'd114, 8'd96, 8'd88, 8'd77, 8'd125, 8'd117, 8'd144, 8'd88, 8'd53, 8'd64, 8'd41, 8'd48, 8'd114, 8'd51, 8'd20, 8'd115, 8'd143, 8'd141, 8'd114, 8'd164, 8'd130, 8'd151, 8'd176, 8'd181, 8'd88, 8'd33, 8'd86, 8'd126, 8'd71, 8'd78, 8'd84, 8'd52, 8'd114, 8'd67, 8'd139, 8'd159, 8'd88, 8'd59, 8'd15, 8'd51, 8'd118, 8'd97, 8'd62, 8'd101, 8'd149, 8'd82, 8'd165, 8'd130, 8'd124, 8'd143, 8'd109, 8'd135, 8'd77, 8'd31, 8'd61, 8'd81, 8'd159, 8'd147, 8'd99, 8'd98, 8'd111, 8'd174, 8'd182, 8'd106, 8'd32, 8'd34, 8'd73, 8'd68, 8'd99, 8'd75, 8'd20, 8'd100, 8'd80, 8'd145, 8'd144, 8'd149, 8'd148, 8'd97, 8'd172, 8'd176, 8'd134, 8'd126, 8'd88, 8'd90, 8'd94, 8'd129, 8'd163, 8'd145, 8'd111, 8'd207, 8'd126, 8'd99, 8'd43, 8'd101, 8'd55, 8'd75, 8'd41, 8'd55, 8'd114, 8'd168, 8'd120, 8'd164, 8'd138, 8'd79, 8'd165, 8'd180, 8'd114, 8'd148, 8'd132, 8'd103, 8'd88, 8'd123, 8'd120, 8'd162, 8'd168, 8'd116, 8'd131, 8'd225, 8'd211, 8'd102, 8'd122, 8'd105, 8'd68, 8'd74, 8'd105, 8'd72, 8'd163, 8'd145, 8'd103, 8'd107, 8'd170, 8'd163, 8'd163, 8'd98, 8'd170, 8'd123, 8'd90, 8'd120, 8'd107, 8'd104, 8'd95, 8'd116, 8'd127, 8'd109, 8'd182, 8'd181, 8'd172, 8'd165, 8'd150, 8'd122, 8'd142, 8'd148, 8'd101, 8'd115, 8'd158, 8'd168, 8'd142, 8'd96, 8'd115, 8'd104, 8'd145, 8'd96, 8'd117, 8'd79, 8'd122, 8'd98, 8'd149, 8'd117, 8'd93, 8'd179, 8'd181, 8'd202, 8'd196, 8'd230, 8'd146, 8'd124, 8'd120, 8'd105, 8'd145, 8'd134, 8'd177, 8'd83, 8'd120, 8'd103, 8'd169, 8'd90, 8'd99, 8'd130, 8'd91, 8'd132, 8'd96, 8'd89, 8'd59, 8'd19, 8'd61, 8'd154, 8'd106, 8'd176, 8'd143, 8'd186, 8'd195, 8'd157, 8'd138, 8'd214, 8'd140, 8'd127, 8'd171, 8'd140, 8'd123, 8'd144, 8'd94, 8'd100, 8'd132, 8'd139, 8'd155, 8'd172, 8'd151, 8'd103, 8'd66, 8'd78, 8'd94, 8'd89, 8'd87, 8'd98, 8'd131, 8'd166, 8'd83, 8'd142, 8'd160, 8'd189, 8'd139, 8'd196, 8'd125, 8'd192, 8'd147, 8'd106, 8'd159, 8'd152, 8'd122, 8'd112, 8'd81, 8'd136, 8'd125, 8'd155, 8'd90, 8'd119, 8'd80, 8'd88, 8'd103, 8'd52, 8'd116, 8'd56, 8'd102, 8'd134, 8'd106, 8'd137, 8'd147, 8'd163, 8'd98, 8'd179, 8'd194, 8'd126, 8'd178, 8'd121, 8'd144, 8'd81, 8'd87, 8'd132, 8'd99, 8'd111, 8'd133, 8'd122, 8'd150, 8'd96, 8'd156, 8'd151, 8'd46, 8'd36, 8'd96, 8'd66, 8'd101, 8'd142, 8'd128, 8'd108, 8'd137, 8'd165, 8'd187, 8'd151, 8'd128, 8'd122, 8'd138, 8'd151, 8'd119, 8'd124, 8'd111, 8'd116, 8'd77, 8'd173, 8'd95, 8'd152, 8'd74, 8'd118, 8'd120, 8'd164, 8'd51, 8'd55, 8'd64, 8'd91, 8'd57, 8'd45, 8'd144, 8'd111, 8'd131, 8'd93, 8'd100, 8'd149, 8'd195, 8'd102, 8'd122, 8'd118, 8'd119, 8'd89, 8'd158, 8'd92, 8'd123, 8'd90, 8'd135, 8'd98, 8'd144, 8'd152, 8'd154, 8'd102, 8'd135, 8'd93, 8'd56, 8'd134, 8'd124, 8'd83, 8'd137, 8'd99, 8'd128, 8'd139, 8'd116, 8'd133, 8'd124, 8'd166, 8'd119, 8'd142, 8'd122, 8'd162, 8'd108, 8'd108, 8'd159, 8'd126, 8'd97, 8'd119, 8'd87, 8'd106, 8'd123, 8'd150, 8'd75, 8'd163, 8'd109, 8'd122, 8'd152, 8'd94, 8'd93, 8'd97, 8'd138, 8'd148, 8'd108, 8'd131, 8'd107, 8'd71, 8'd79, 8'd141, 8'd94, 8'd97, 8'd95, 8'd141, 8'd117, 8'd126, 8'd150, 8'd146, 8'd164, 8'd78, 8'd118, 8'd95, 8'd80, 8'd154, 8'd85, 8'd87, 8'd91, 8'd124, 8'd84, 8'd157, 8'd149, 8'd170, 8'd154, 8'd170, 8'd96, 8'd92, 8'd125, 8'd115, 8'd167, 8'd143, 8'd108, 8'd108, 8'd83, 8'd83, 8'd123, 8'd95, 8'd121})
) cell_0_50 (
    .clk(clk),
    .input_index(index_0_49_50),
    .input_value(value_0_49_50),
    .input_result(result_0_49_50),
    .input_enable(enable_0_49_50),
    .output_index(index_0_50_51),
    .output_value(value_0_50_51),
    .output_result(result_0_50_51),
    .output_enable(enable_0_50_51)
);

wire [10-1:0] index_0_51_52;
wire [`DATA_WIDTH-1:0] value_0_51_52;
wire [`DATA_WIDTH*4:0] result_0_51_52;
wire enable_0_51_52;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd147, 8'd129, 8'd155, 8'd162, 8'd148, 8'd135, 8'd112, 8'd106, 8'd69, 8'd73, 8'd72, 8'd96, 8'd111, 8'd120, 8'd108, 8'd67, 8'd122, 8'd102, 8'd103, 8'd108, 8'd131, 8'd99, 8'd81, 8'd102, 8'd121, 8'd98, 8'd104, 8'd108, 8'd75, 8'd79, 8'd106, 8'd149, 8'd167, 8'd154, 8'd144, 8'd80, 8'd91, 8'd129, 8'd86, 8'd76, 8'd80, 8'd95, 8'd169, 8'd154, 8'd85, 8'd142, 8'd92, 8'd156, 8'd113, 8'd174, 8'd115, 8'd102, 8'd167, 8'd133, 8'd140, 8'd128, 8'd87, 8'd132, 8'd173, 8'd79, 8'd95, 8'd172, 8'd137, 8'd175, 8'd141, 8'd102, 8'd91, 8'd97, 8'd95, 8'd69, 8'd155, 8'd108, 8'd68, 8'd96, 8'd67, 8'd154, 8'd140, 8'd152, 8'd158, 8'd152, 8'd130, 8'd155, 8'd105, 8'd134, 8'd98, 8'd105, 8'd158, 8'd168, 8'd111, 8'd178, 8'd87, 8'd107, 8'd71, 8'd124, 8'd147, 8'd145, 8'd117, 8'd101, 8'd128, 8'd143, 8'd164, 8'd97, 8'd82, 8'd139, 8'd107, 8'd34, 8'd60, 8'd62, 8'd55, 8'd90, 8'd109, 8'd87, 8'd168, 8'd106, 8'd89, 8'd135, 8'd190, 8'd182, 8'd118, 8'd149, 8'd141, 8'd108, 8'd148, 8'd100, 8'd138, 8'd162, 8'd186, 8'd184, 8'd178, 8'd173, 8'd165, 8'd123, 8'd102, 8'd98, 8'd111, 8'd83, 8'd128, 8'd110, 8'd146, 8'd146, 8'd143, 8'd86, 8'd170, 8'd113, 8'd99, 8'd106, 8'd79, 8'd155, 8'd91, 8'd99, 8'd153, 8'd110, 8'd158, 8'd152, 8'd161, 8'd177, 8'd183, 8'd170, 8'd100, 8'd144, 8'd144, 8'd153, 8'd65, 8'd136, 8'd98, 8'd126, 8'd85, 8'd108, 8'd160, 8'd137, 8'd168, 8'd89, 8'd170, 8'd136, 8'd126, 8'd79, 8'd94, 8'd86, 8'd113, 8'd95, 8'd128, 8'd169, 8'd88, 8'd187, 8'd129, 8'd151, 8'd165, 8'd94, 8'd134, 8'd123, 8'd128, 8'd143, 8'd142, 8'd92, 8'd94, 8'd127, 8'd136, 8'd162, 8'd168, 8'd154, 8'd148, 8'd155, 8'd137, 8'd142, 8'd97, 8'd86, 8'd146, 8'd114, 8'd95, 8'd88, 8'd88, 8'd92, 8'd134, 8'd147, 8'd100, 8'd116, 8'd128, 8'd121, 8'd100, 8'd171, 8'd65, 8'd101, 8'd96, 8'd128, 8'd82, 8'd162, 8'd139, 8'd153, 8'd180, 8'd175, 8'd95, 8'd153, 8'd86, 8'd145, 8'd81, 8'd124, 8'd154, 8'd96, 8'd71, 8'd108, 8'd141, 8'd129, 8'd150, 8'd116, 8'd135, 8'd132, 8'd94, 8'd89, 8'd51, 8'd71, 8'd116, 8'd149, 8'd81, 8'd83, 8'd103, 8'd176, 8'd159, 8'd123, 8'd90, 8'd98, 8'd97, 8'd93, 8'd118, 8'd160, 8'd125, 8'd123, 8'd52, 8'd78, 8'd158, 8'd193, 8'd170, 8'd164, 8'd90, 8'd136, 8'd147, 8'd106, 8'd114, 8'd90, 8'd77, 8'd115, 8'd141, 8'd151, 8'd190, 8'd189, 8'd122, 8'd167, 8'd151, 8'd164, 8'd84, 8'd122, 8'd127, 8'd138, 8'd97, 8'd64, 8'd123, 8'd104, 8'd147, 8'd161, 8'd137, 8'd116, 8'd144, 8'd114, 8'd141, 8'd78, 8'd116, 8'd153, 8'd133, 8'd141, 8'd116, 8'd161, 8'd161, 8'd128, 8'd138, 8'd145, 8'd159, 8'd163, 8'd151, 8'd130, 8'd94, 8'd108, 8'd115, 8'd97, 8'd73, 8'd103, 8'd195, 8'd107, 8'd152, 8'd92, 8'd154, 8'd83, 8'd135, 8'd153, 8'd150, 8'd87, 8'd95, 8'd117, 8'd140, 8'd106, 8'd126, 8'd106, 8'd143, 8'd141, 8'd96, 8'd88, 8'd112, 8'd118, 8'd112, 8'd138, 8'd142, 8'd46, 8'd148, 8'd102, 8'd123, 8'd125, 8'd125, 8'd113, 8'd110, 8'd165, 8'd93, 8'd65, 8'd103, 8'd118, 8'd97, 8'd144, 8'd152, 8'd170, 8'd123, 8'd128, 8'd96, 8'd121, 8'd106, 8'd164, 8'd69, 8'd122, 8'd112, 8'd135, 8'd135, 8'd111, 8'd131, 8'd155, 8'd111, 8'd104, 8'd127, 8'd167, 8'd107, 8'd125, 8'd78, 8'd127, 8'd144, 8'd105, 8'd92, 8'd128, 8'd132, 8'd110, 8'd121, 8'd184, 8'd144, 8'd171, 8'd85, 8'd131, 8'd121, 8'd157, 8'd74, 8'd63, 8'd50, 8'd60, 8'd102, 8'd84, 8'd123, 8'd158, 8'd88, 8'd108, 8'd127, 8'd127, 8'd138, 8'd69, 8'd126, 8'd126, 8'd109, 8'd131, 8'd147, 8'd136, 8'd129, 8'd126, 8'd133, 8'd132, 8'd147, 8'd90, 8'd104, 8'd127, 8'd88, 8'd102, 8'd46, 8'd96, 8'd143, 8'd147, 8'd152, 8'd159, 8'd71, 8'd98, 8'd86, 8'd78, 8'd161, 8'd136, 8'd58, 8'd79, 8'd87, 8'd103, 8'd69, 8'd67, 8'd69, 8'd110, 8'd149, 8'd99, 8'd120, 8'd167, 8'd175, 8'd162, 8'd109, 8'd34, 8'd78, 8'd139, 8'd112, 8'd116, 8'd130, 8'd85, 8'd125, 8'd79, 8'd156, 8'd85, 8'd92, 8'd121, 8'd50, 8'd131, 8'd128, 8'd117, 8'd121, 8'd95, 8'd76, 8'd167, 8'd135, 8'd107, 8'd152, 8'd160, 8'd124, 8'd168, 8'd145, 8'd134, 8'd97, 8'd130, 8'd108, 8'd159, 8'd88, 8'd142, 8'd131, 8'd74, 8'd92, 8'd86, 8'd88, 8'd102, 8'd138, 8'd103, 8'd66, 8'd137, 8'd68, 8'd106, 8'd141, 8'd157, 8'd192, 8'd174, 8'd79, 8'd133, 8'd121, 8'd103, 8'd116, 8'd70, 8'd117, 8'd129, 8'd117, 8'd137, 8'd154, 8'd138, 8'd103, 8'd83, 8'd152, 8'd86, 8'd87, 8'd97, 8'd141, 8'd120, 8'd76, 8'd87, 8'd144, 8'd163, 8'd83, 8'd146, 8'd144, 8'd128, 8'd170, 8'd152, 8'd126, 8'd125, 8'd109, 8'd134, 8'd142, 8'd162, 8'd173, 8'd106, 8'd156, 8'd159, 8'd92, 8'd156, 8'd98, 8'd151, 8'd118, 8'd100, 8'd77, 8'd112, 8'd148, 8'd94, 8'd115, 8'd82, 8'd83, 8'd166, 8'd113, 8'd77, 8'd138, 8'd151, 8'd75, 8'd176, 8'd146, 8'd115, 8'd163, 8'd128, 8'd167, 8'd143, 8'd120, 8'd85, 8'd103, 8'd142, 8'd118, 8'd84, 8'd60, 8'd122, 8'd136, 8'd151, 8'd147, 8'd75, 8'd81, 8'd94, 8'd152, 8'd91, 8'd149, 8'd105, 8'd100, 8'd89, 8'd85, 8'd168, 8'd118, 8'd171, 8'd149, 8'd128, 8'd103, 8'd167, 8'd129, 8'd93, 8'd146, 8'd158, 8'd82, 8'd137, 8'd113, 8'd111, 8'd147, 8'd83, 8'd143, 8'd117, 8'd164, 8'd162, 8'd90, 8'd126, 8'd57, 8'd93, 8'd157, 8'd155, 8'd136, 8'd110, 8'd118, 8'd179, 8'd134, 8'd98, 8'd114, 8'd109, 8'd99, 8'd169, 8'd151, 8'd81, 8'd113, 8'd56, 8'd52, 8'd114, 8'd129, 8'd99, 8'd122, 8'd105, 8'd110, 8'd94, 8'd164, 8'd123, 8'd100, 8'd84, 8'd97, 8'd135, 8'd88, 8'd87, 8'd147, 8'd135, 8'd89, 8'd143, 8'd129, 8'd108, 8'd151, 8'd161, 8'd147, 8'd151, 8'd90, 8'd97, 8'd109, 8'd68, 8'd68, 8'd82, 8'd150, 8'd112, 8'd122, 8'd105, 8'd135, 8'd152, 8'd178, 8'd123, 8'd94, 8'd108, 8'd145, 8'd80, 8'd118, 8'd90, 8'd164, 8'd118, 8'd165, 8'd185, 8'd158, 8'd150, 8'd197, 8'd118, 8'd100, 8'd76, 8'd138, 8'd137, 8'd93, 8'd81, 8'd101, 8'd72, 8'd162, 8'd123, 8'd174, 8'd123, 8'd146, 8'd123, 8'd184, 8'd136, 8'd96, 8'd156, 8'd125, 8'd114, 8'd133, 8'd181, 8'd155, 8'd151, 8'd158, 8'd198, 8'd154, 8'd183, 8'd117, 8'd183, 8'd110, 8'd101, 8'd88, 8'd95, 8'd122, 8'd97, 8'd82, 8'd85, 8'd135, 8'd76, 8'd92, 8'd163, 8'd158, 8'd159, 8'd159, 8'd98, 8'd155, 8'd104, 8'd171, 8'd122, 8'd179, 8'd119, 8'd186, 8'd180, 8'd100, 8'd157, 8'd97, 8'd97, 8'd122, 8'd94, 8'd169, 8'd135, 8'd75, 8'd134, 8'd82, 8'd104, 8'd105, 8'd160, 8'd165, 8'd141, 8'd102, 8'd71, 8'd115, 8'd108, 8'd147, 8'd138, 8'd106, 8'd108, 8'd134, 8'd120, 8'd88, 8'd91, 8'd135, 8'd120, 8'd100, 8'd96, 8'd170, 8'd104, 8'd169, 8'd156, 8'd81, 8'd120})
) cell_0_51 (
    .clk(clk),
    .input_index(index_0_50_51),
    .input_value(value_0_50_51),
    .input_result(result_0_50_51),
    .input_enable(enable_0_50_51),
    .output_index(index_0_51_52),
    .output_value(value_0_51_52),
    .output_result(result_0_51_52),
    .output_enable(enable_0_51_52)
);

wire [10-1:0] index_0_52_53;
wire [`DATA_WIDTH-1:0] value_0_52_53;
wire [`DATA_WIDTH*4:0] result_0_52_53;
wire enable_0_52_53;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd159, 8'd108, 8'd104, 8'd84, 8'd157, 8'd88, 8'd111, 8'd159, 8'd154, 8'd196, 8'd186, 8'd151, 8'd201, 8'd161, 8'd193, 8'd144, 8'd152, 8'd164, 8'd97, 8'd186, 8'd177, 8'd94, 8'd121, 8'd171, 8'd85, 8'd106, 8'd128, 8'd117, 8'd96, 8'd125, 8'd156, 8'd101, 8'd107, 8'd162, 8'd168, 8'd111, 8'd98, 8'd146, 8'd146, 8'd176, 8'd144, 8'd176, 8'd113, 8'd125, 8'd127, 8'd162, 8'd156, 8'd182, 8'd104, 8'd140, 8'd172, 8'd113, 8'd162, 8'd152, 8'd148, 8'd86, 8'd75, 8'd153, 8'd124, 8'd126, 8'd64, 8'd74, 8'd81, 8'd109, 8'd101, 8'd132, 8'd78, 8'd140, 8'd90, 8'd148, 8'd109, 8'd176, 8'd111, 8'd148, 8'd121, 8'd112, 8'd114, 8'd168, 8'd108, 8'd78, 8'd107, 8'd150, 8'd93, 8'd105, 8'd75, 8'd158, 8'd106, 8'd139, 8'd132, 8'd154, 8'd130, 8'd101, 8'd102, 8'd116, 8'd118, 8'd149, 8'd140, 8'd82, 8'd168, 8'd153, 8'd163, 8'd99, 8'd152, 8'd164, 8'd115, 8'd158, 8'd146, 8'd65, 8'd100, 8'd124, 8'd84, 8'd98, 8'd127, 8'd146, 8'd150, 8'd163, 8'd135, 8'd162, 8'd133, 8'd94, 8'd137, 8'd114, 8'd116, 8'd98, 8'd100, 8'd71, 8'd122, 8'd101, 8'd116, 8'd125, 8'd80, 8'd76, 8'd161, 8'd161, 8'd124, 8'd81, 8'd81, 8'd99, 8'd82, 8'd97, 8'd71, 8'd93, 8'd151, 8'd122, 8'd131, 8'd111, 8'd178, 8'd111, 8'd78, 8'd103, 8'd80, 8'd133, 8'd98, 8'd90, 8'd108, 8'd120, 8'd154, 8'd140, 8'd81, 8'd164, 8'd178, 8'd95, 8'd92, 8'd154, 8'd154, 8'd123, 8'd152, 8'd81, 8'd130, 8'd85, 8'd87, 8'd128, 8'd118, 8'd91, 8'd118, 8'd136, 8'd92, 8'd83, 8'd85, 8'd114, 8'd146, 8'd95, 8'd80, 8'd129, 8'd138, 8'd156, 8'd116, 8'd89, 8'd136, 8'd96, 8'd134, 8'd81, 8'd118, 8'd124, 8'd122, 8'd86, 8'd162, 8'd113, 8'd145, 8'd164, 8'd135, 8'd143, 8'd85, 8'd157, 8'd152, 8'd94, 8'd156, 8'd84, 8'd117, 8'd97, 8'd164, 8'd155, 8'd61, 8'd99, 8'd66, 8'd93, 8'd118, 8'd146, 8'd146, 8'd142, 8'd63, 8'd71, 8'd89, 8'd149, 8'd179, 8'd125, 8'd125, 8'd118, 8'd123, 8'd125, 8'd137, 8'd157, 8'd115, 8'd105, 8'd82, 8'd149, 8'd146, 8'd152, 8'd97, 8'd94, 8'd131, 8'd138, 8'd137, 8'd63, 8'd81, 8'd129, 8'd86, 8'd134, 8'd131, 8'd89, 8'd114, 8'd154, 8'd89, 8'd121, 8'd123, 8'd111, 8'd104, 8'd118, 8'd133, 8'd144, 8'd90, 8'd112, 8'd87, 8'd89, 8'd178, 8'd158, 8'd185, 8'd192, 8'd152, 8'd78, 8'd129, 8'd157, 8'd66, 8'd61, 8'd121, 8'd130, 8'd136, 8'd119, 8'd88, 8'd166, 8'd124, 8'd175, 8'd162, 8'd96, 8'd137, 8'd157, 8'd122, 8'd75, 8'd152, 8'd136, 8'd120, 8'd117, 8'd111, 8'd118, 8'd151, 8'd208, 8'd108, 8'd92, 8'd80, 8'd98, 8'd141, 8'd84, 8'd86, 8'd170, 8'd168, 8'd158, 8'd74, 8'd82, 8'd150, 8'd217, 8'd171, 8'd93, 8'd71, 8'd127, 8'd153, 8'd147, 8'd121, 8'd116, 8'd146, 8'd144, 8'd147, 8'd158, 8'd189, 8'd157, 8'd98, 8'd146, 8'd97, 8'd150, 8'd129, 8'd144, 8'd94, 8'd117, 8'd97, 8'd97, 8'd64, 8'd98, 8'd88, 8'd166, 8'd163, 8'd129, 8'd138, 8'd79, 8'd84, 8'd108, 8'd122, 8'd136, 8'd165, 8'd154, 8'd147, 8'd169, 8'd130, 8'd112, 8'd93, 8'd64, 8'd132, 8'd134, 8'd129, 8'd138, 8'd132, 8'd108, 8'd146, 8'd151, 8'd98, 8'd79, 8'd165, 8'd182, 8'd114, 8'd115, 8'd76, 8'd135, 8'd155, 8'd131, 8'd132, 8'd115, 8'd122, 8'd112, 8'd119, 8'd193, 8'd126, 8'd138, 8'd117, 8'd72, 8'd61, 8'd121, 8'd80, 8'd58, 8'd123, 8'd99, 8'd188, 8'd184, 8'd101, 8'd154, 8'd148, 8'd190, 8'd184, 8'd137, 8'd71, 8'd128, 8'd118, 8'd100, 8'd101, 8'd175, 8'd165, 8'd192, 8'd193, 8'd93, 8'd125, 8'd65, 8'd42, 8'd107, 8'd53, 8'd103, 8'd55, 8'd96, 8'd142, 8'd165, 8'd188, 8'd98, 8'd171, 8'd174, 8'd105, 8'd133, 8'd178, 8'd96, 8'd95, 8'd144, 8'd148, 8'd108, 8'd125, 8'd145, 8'd174, 8'd182, 8'd153, 8'd161, 8'd108, 8'd80, 8'd59, 8'd55, 8'd103, 8'd76, 8'd138, 8'd97, 8'd142, 8'd126, 8'd153, 8'd136, 8'd101, 8'd122, 8'd110, 8'd60, 8'd41, 8'd128, 8'd136, 8'd130, 8'd153, 8'd141, 8'd124, 8'd96, 8'd102, 8'd128, 8'd112, 8'd136, 8'd77, 8'd137, 8'd107, 8'd156, 8'd110, 8'd82, 8'd145, 8'd110, 8'd132, 8'd135, 8'd150, 8'd118, 8'd83, 8'd163, 8'd164, 8'd47, 8'd72, 8'd17, 8'd129, 8'd156, 8'd129, 8'd100, 8'd149, 8'd188, 8'd165, 8'd119, 8'd104, 8'd71, 8'd131, 8'd117, 8'd156, 8'd110, 8'd113, 8'd163, 8'd82, 8'd181, 8'd136, 8'd162, 8'd188, 8'd120, 8'd126, 8'd145, 8'd78, 8'd108, 8'd106, 8'd71, 8'd117, 8'd134, 8'd101, 8'd144, 8'd170, 8'd147, 8'd135, 8'd130, 8'd170, 8'd161, 8'd135, 8'd139, 8'd131, 8'd163, 8'd100, 8'd138, 8'd120, 8'd168, 8'd183, 8'd175, 8'd141, 8'd157, 8'd109, 8'd149, 8'd152, 8'd89, 8'd68, 8'd125, 8'd67, 8'd80, 8'd92, 8'd77, 8'd91, 8'd139, 8'd131, 8'd138, 8'd91, 8'd140, 8'd165, 8'd169, 8'd168, 8'd116, 8'd136, 8'd110, 8'd185, 8'd144, 8'd178, 8'd116, 8'd151, 8'd92, 8'd144, 8'd155, 8'd141, 8'd76, 8'd88, 8'd132, 8'd140, 8'd112, 8'd102, 8'd83, 8'd85, 8'd109, 8'd118, 8'd157, 8'd107, 8'd75, 8'd127, 8'd175, 8'd114, 8'd104, 8'd115, 8'd192, 8'd181, 8'd171, 8'd104, 8'd195, 8'd195, 8'd116, 8'd74, 8'd75, 8'd116, 8'd96, 8'd83, 8'd121, 8'd68, 8'd89, 8'd124, 8'd98, 8'd100, 8'd156, 8'd67, 8'd124, 8'd120, 8'd163, 8'd86, 8'd91, 8'd153, 8'd93, 8'd99, 8'd95, 8'd91, 8'd94, 8'd143, 8'd156, 8'd130, 8'd113, 8'd161, 8'd132, 8'd81, 8'd105, 8'd149, 8'd103, 8'd119, 8'd136, 8'd114, 8'd115, 8'd61, 8'd104, 8'd87, 8'd104, 8'd82, 8'd81, 8'd128, 8'd105, 8'd163, 8'd111, 8'd170, 8'd162, 8'd169, 8'd99, 8'd134, 8'd129, 8'd117, 8'd78, 8'd152, 8'd117, 8'd122, 8'd139, 8'd65, 8'd70, 8'd79, 8'd111, 8'd105, 8'd118, 8'd111, 8'd116, 8'd77, 8'd132, 8'd101, 8'd105, 8'd125, 8'd77, 8'd113, 8'd168, 8'd137, 8'd167, 8'd170, 8'd156, 8'd98, 8'd138, 8'd165, 8'd122, 8'd69, 8'd163, 8'd135, 8'd95, 8'd100, 8'd102, 8'd73, 8'd141, 8'd109, 8'd70, 8'd123, 8'd81, 8'd66, 8'd139, 8'd134, 8'd140, 8'd116, 8'd82, 8'd119, 8'd146, 8'd132, 8'd118, 8'd89, 8'd87, 8'd128, 8'd114, 8'd117, 8'd138, 8'd76, 8'd114, 8'd143, 8'd90, 8'd74, 8'd98, 8'd125, 8'd97, 8'd95, 8'd145, 8'd110, 8'd152, 8'd129, 8'd129, 8'd121, 8'd130, 8'd79, 8'd142, 8'd93, 8'd79, 8'd69, 8'd127, 8'd106, 8'd67, 8'd99, 8'd98, 8'd73, 8'd123, 8'd79, 8'd75, 8'd125, 8'd89, 8'd106, 8'd98, 8'd119, 8'd140, 8'd66, 8'd73, 8'd57, 8'd89, 8'd78, 8'd169, 8'd129, 8'd151, 8'd100, 8'd115, 8'd137, 8'd106, 8'd104, 8'd121, 8'd144, 8'd113, 8'd65, 8'd79, 8'd119, 8'd126, 8'd167, 8'd137, 8'd169, 8'd105, 8'd140, 8'd79, 8'd133, 8'd73, 8'd81, 8'd79, 8'd115, 8'd121, 8'd93, 8'd158, 8'd82, 8'd122, 8'd86, 8'd138, 8'd75, 8'd120, 8'd74, 8'd83, 8'd134, 8'd103, 8'd82, 8'd80, 8'd101, 8'd166, 8'd127, 8'd81})
) cell_0_52 (
    .clk(clk),
    .input_index(index_0_51_52),
    .input_value(value_0_51_52),
    .input_result(result_0_51_52),
    .input_enable(enable_0_51_52),
    .output_index(index_0_52_53),
    .output_value(value_0_52_53),
    .output_result(result_0_52_53),
    .output_enable(enable_0_52_53)
);

wire [10-1:0] index_0_53_54;
wire [`DATA_WIDTH-1:0] value_0_53_54;
wire [`DATA_WIDTH*4:0] result_0_53_54;
wire enable_0_53_54;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd111, 8'd161, 8'd77, 8'd143, 8'd105, 8'd154, 8'd146, 8'd149, 8'd81, 8'd98, 8'd107, 8'd144, 8'd133, 8'd98, 8'd90, 8'd144, 8'd119, 8'd152, 8'd133, 8'd102, 8'd89, 8'd84, 8'd147, 8'd144, 8'd149, 8'd109, 8'd103, 8'd110, 8'd76, 8'd160, 8'd124, 8'd92, 8'd96, 8'd100, 8'd110, 8'd71, 8'd141, 8'd120, 8'd90, 8'd79, 8'd131, 8'd89, 8'd124, 8'd65, 8'd113, 8'd90, 8'd99, 8'd61, 8'd75, 8'd101, 8'd132, 8'd86, 8'd122, 8'd132, 8'd117, 8'd131, 8'd166, 8'd107, 8'd173, 8'd153, 8'd168, 8'd147, 8'd95, 8'd136, 8'd127, 8'd146, 8'd95, 8'd149, 8'd121, 8'd119, 8'd129, 8'd162, 8'd127, 8'd132, 8'd92, 8'd168, 8'd105, 8'd108, 8'd96, 8'd99, 8'd143, 8'd76, 8'd156, 8'd136, 8'd90, 8'd140, 8'd112, 8'd109, 8'd99, 8'd140, 8'd164, 8'd152, 8'd155, 8'd101, 8'd122, 8'd169, 8'd180, 8'd116, 8'd173, 8'd136, 8'd166, 8'd153, 8'd101, 8'd160, 8'd141, 8'd153, 8'd126, 8'd152, 8'd131, 8'd118, 8'd74, 8'd109, 8'd83, 8'd170, 8'd94, 8'd88, 8'd151, 8'd90, 8'd144, 8'd151, 8'd166, 8'd158, 8'd145, 8'd98, 8'd82, 8'd95, 8'd117, 8'd106, 8'd93, 8'd119, 8'd98, 8'd170, 8'd166, 8'd129, 8'd169, 8'd135, 8'd200, 8'd86, 8'd132, 8'd76, 8'd165, 8'd168, 8'd99, 8'd111, 8'd162, 8'd134, 8'd92, 8'd180, 8'd121, 8'd98, 8'd159, 8'd118, 8'd115, 8'd136, 8'd161, 8'd151, 8'd90, 8'd89, 8'd158, 8'd140, 8'd115, 8'd147, 8'd77, 8'd126, 8'd170, 8'd112, 8'd118, 8'd74, 8'd77, 8'd136, 8'd162, 8'd121, 8'd162, 8'd84, 8'd157, 8'd164, 8'd101, 8'd156, 8'd164, 8'd132, 8'd80, 8'd167, 8'd110, 8'd80, 8'd159, 8'd121, 8'd101, 8'd162, 8'd96, 8'd113, 8'd161, 8'd153, 8'd132, 8'd101, 8'd128, 8'd85, 8'd162, 8'd157, 8'd149, 8'd137, 8'd138, 8'd99, 8'd160, 8'd173, 8'd127, 8'd174, 8'd140, 8'd145, 8'd115, 8'd83, 8'd158, 8'd111, 8'd133, 8'd91, 8'd136, 8'd175, 8'd93, 8'd188, 8'd130, 8'd167, 8'd127, 8'd184, 8'd157, 8'd88, 8'd157, 8'd185, 8'd150, 8'd114, 8'd151, 8'd168, 8'd112, 8'd122, 8'd179, 8'd92, 8'd144, 8'd156, 8'd142, 8'd174, 8'd111, 8'd110, 8'd156, 8'd122, 8'd93, 8'd143, 8'd117, 8'd188, 8'd104, 8'd167, 8'd119, 8'd138, 8'd131, 8'd124, 8'd109, 8'd125, 8'd174, 8'd179, 8'd130, 8'd127, 8'd142, 8'd91, 8'd96, 8'd126, 8'd179, 8'd115, 8'd94, 8'd80, 8'd129, 8'd78, 8'd136, 8'd126, 8'd127, 8'd128, 8'd138, 8'd151, 8'd144, 8'd157, 8'd217, 8'd106, 8'd107, 8'd118, 8'd139, 8'd164, 8'd163, 8'd159, 8'd172, 8'd155, 8'd159, 8'd153, 8'd90, 8'd146, 8'd95, 8'd125, 8'd96, 8'd60, 8'd140, 8'd142, 8'd141, 8'd124, 8'd72, 8'd95, 8'd90, 8'd154, 8'd115, 8'd174, 8'd149, 8'd111, 8'd100, 8'd73, 8'd150, 8'd174, 8'd146, 8'd201, 8'd128, 8'd107, 8'd167, 8'd101, 8'd182, 8'd116, 8'd93, 8'd72, 8'd115, 8'd140, 8'd91, 8'd125, 8'd113, 8'd129, 8'd71, 8'd98, 8'd121, 8'd112, 8'd110, 8'd148, 8'd187, 8'd125, 8'd79, 8'd98, 8'd179, 8'd110, 8'd95, 8'd149, 8'd177, 8'd155, 8'd129, 8'd80, 8'd112, 8'd160, 8'd148, 8'd146, 8'd130, 8'd122, 8'd74, 8'd104, 8'd147, 8'd151, 8'd132, 8'd148, 8'd143, 8'd105, 8'd138, 8'd89, 8'd146, 8'd174, 8'd164, 8'd121, 8'd83, 8'd148, 8'd161, 8'd144, 8'd103, 8'd106, 8'd93, 8'd79, 8'd131, 8'd157, 8'd88, 8'd99, 8'd156, 8'd102, 8'd166, 8'd167, 8'd99, 8'd91, 8'd125, 8'd107, 8'd89, 8'd52, 8'd122, 8'd128, 8'd150, 8'd118, 8'd101, 8'd112, 8'd156, 8'd185, 8'd161, 8'd117, 8'd124, 8'd58, 8'd70, 8'd98, 8'd100, 8'd130, 8'd87, 8'd87, 8'd82, 8'd131, 8'd103, 8'd72, 8'd116, 8'd121, 8'd127, 8'd109, 8'd132, 8'd116, 8'd107, 8'd64, 8'd93, 8'd123, 8'd150, 8'd115, 8'd111, 8'd137, 8'd100, 8'd73, 8'd11, 8'd47, 8'd39, 8'd103, 8'd96, 8'd88, 8'd72, 8'd131, 8'd64, 8'd100, 8'd66, 8'd89, 8'd89, 8'd130, 8'd117, 8'd132, 8'd129, 8'd91, 8'd55, 8'd87, 8'd85, 8'd160, 8'd150, 8'd115, 8'd153, 8'd129, 8'd197, 8'd117, 8'd112, 8'd38, 8'd65, 8'd86, 8'd85, 8'd119, 8'd82, 8'd109, 8'd153, 8'd86, 8'd124, 8'd107, 8'd139, 8'd133, 8'd92, 8'd118, 8'd123, 8'd127, 8'd90, 8'd113, 8'd179, 8'd86, 8'd157, 8'd115, 8'd174, 8'd115, 8'd213, 8'd188, 8'd152, 8'd76, 8'd100, 8'd105, 8'd78, 8'd169, 8'd84, 8'd97, 8'd166, 8'd70, 8'd150, 8'd92, 8'd150, 8'd103, 8'd155, 8'd112, 8'd101, 8'd142, 8'd83, 8'd140, 8'd157, 8'd153, 8'd91, 8'd166, 8'd143, 8'd184, 8'd147, 8'd108, 8'd126, 8'd99, 8'd122, 8'd128, 8'd156, 8'd135, 8'd115, 8'd141, 8'd137, 8'd146, 8'd145, 8'd165, 8'd113, 8'd121, 8'd99, 8'd110, 8'd153, 8'd100, 8'd143, 8'd115, 8'd92, 8'd93, 8'd103, 8'd101, 8'd165, 8'd91, 8'd115, 8'd153, 8'd119, 8'd149, 8'd150, 8'd141, 8'd123, 8'd161, 8'd173, 8'd105, 8'd148, 8'd129, 8'd160, 8'd101, 8'd102, 8'd176, 8'd128, 8'd142, 8'd120, 8'd87, 8'd139, 8'd150, 8'd182, 8'd76, 8'd93, 8'd127, 8'd107, 8'd115, 8'd157, 8'd126, 8'd108, 8'd157, 8'd105, 8'd121, 8'd153, 8'd99, 8'd163, 8'd107, 8'd147, 8'd150, 8'd111, 8'd177, 8'd118, 8'd92, 8'd162, 8'd87, 8'd162, 8'd104, 8'd168, 8'd92, 8'd117, 8'd79, 8'd181, 8'd90, 8'd149, 8'd100, 8'd90, 8'd152, 8'd102, 8'd84, 8'd153, 8'd110, 8'd154, 8'd167, 8'd96, 8'd115, 8'd156, 8'd166, 8'd91, 8'd140, 8'd110, 8'd91, 8'd127, 8'd176, 8'd94, 8'd151, 8'd155, 8'd132, 8'd132, 8'd148, 8'd165, 8'd81, 8'd140, 8'd144, 8'd176, 8'd145, 8'd121, 8'd136, 8'd81, 8'd84, 8'd98, 8'd166, 8'd138, 8'd118, 8'd147, 8'd142, 8'd163, 8'd107, 8'd89, 8'd124, 8'd139, 8'd99, 8'd174, 8'd87, 8'd178, 8'd137, 8'd141, 8'd141, 8'd91, 8'd90, 8'd67, 8'd76, 8'd94, 8'd155, 8'd137, 8'd130, 8'd79, 8'd74, 8'd143, 8'd169, 8'd144, 8'd168, 8'd179, 8'd129, 8'd106, 8'd105, 8'd124, 8'd136, 8'd136, 8'd164, 8'd96, 8'd130, 8'd81, 8'd151, 8'd150, 8'd112, 8'd125, 8'd162, 8'd72, 8'd133, 8'd153, 8'd81, 8'd123, 8'd136, 8'd120, 8'd101, 8'd152, 8'd178, 8'd124, 8'd155, 8'd167, 8'd181, 8'd196, 8'd116, 8'd127, 8'd119, 8'd86, 8'd101, 8'd84, 8'd107, 8'd133, 8'd71, 8'd103, 8'd67, 8'd167, 8'd120, 8'd124, 8'd95, 8'd118, 8'd150, 8'd81, 8'd135, 8'd135, 8'd108, 8'd79, 8'd144, 8'd110, 8'd153, 8'd110, 8'd67, 8'd77, 8'd121, 8'd143, 8'd61, 8'd124, 8'd89, 8'd121, 8'd143, 8'd153, 8'd119, 8'd91, 8'd116, 8'd145, 8'd128, 8'd104, 8'd144, 8'd72, 8'd70, 8'd62, 8'd108, 8'd150, 8'd70, 8'd117, 8'd92, 8'd150, 8'd160, 8'd93, 8'd69, 8'd120, 8'd92, 8'd120, 8'd137, 8'd60, 8'd98, 8'd144, 8'd122, 8'd71, 8'd140, 8'd163, 8'd129, 8'd87, 8'd117, 8'd115, 8'd101, 8'd146, 8'd158, 8'd117, 8'd130, 8'd155, 8'd103, 8'd118, 8'd158, 8'd113, 8'd134, 8'd93, 8'd153, 8'd140, 8'd114, 8'd124, 8'd129, 8'd82, 8'd164, 8'd108, 8'd106, 8'd101, 8'd127, 8'd106, 8'd76, 8'd139, 8'd107})
) cell_0_53 (
    .clk(clk),
    .input_index(index_0_52_53),
    .input_value(value_0_52_53),
    .input_result(result_0_52_53),
    .input_enable(enable_0_52_53),
    .output_index(index_0_53_54),
    .output_value(value_0_53_54),
    .output_result(result_0_53_54),
    .output_enable(enable_0_53_54)
);

wire [10-1:0] index_0_54_55;
wire [`DATA_WIDTH-1:0] value_0_54_55;
wire [`DATA_WIDTH*4:0] result_0_54_55;
wire enable_0_54_55;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd116, 8'd156, 8'd117, 8'd146, 8'd154, 8'd111, 8'd163, 8'd155, 8'd150, 8'd93, 8'd138, 8'd150, 8'd159, 8'd104, 8'd162, 8'd92, 8'd115, 8'd88, 8'd134, 8'd154, 8'd128, 8'd155, 8'd79, 8'd86, 8'd119, 8'd144, 8'd125, 8'd155, 8'd169, 8'd119, 8'd125, 8'd103, 8'd80, 8'd91, 8'd112, 8'd101, 8'd149, 8'd125, 8'd95, 8'd111, 8'd94, 8'd151, 8'd127, 8'd111, 8'd90, 8'd109, 8'd153, 8'd158, 8'd119, 8'd148, 8'd109, 8'd151, 8'd154, 8'd149, 8'd88, 8'd97, 8'd75, 8'd73, 8'd110, 8'd77, 8'd59, 8'd100, 8'd70, 8'd108, 8'd106, 8'd61, 8'd79, 8'd110, 8'd135, 8'd127, 8'd117, 8'd105, 8'd157, 8'd116, 8'd205, 8'd187, 8'd181, 8'd158, 8'd127, 8'd140, 8'd173, 8'd106, 8'd165, 8'd133, 8'd147, 8'd120, 8'd79, 8'd83, 8'd78, 8'd117, 8'd128, 8'd150, 8'd144, 8'd154, 8'd118, 8'd93, 8'd117, 8'd124, 8'd162, 8'd85, 8'd151, 8'd176, 8'd114, 8'd121, 8'd196, 8'd218, 8'd138, 8'd121, 8'd108, 8'd102, 8'd110, 8'd100, 8'd102, 8'd153, 8'd88, 8'd66, 8'd82, 8'd93, 8'd111, 8'd97, 8'd148, 8'd152, 8'd127, 8'd168, 8'd68, 8'd90, 8'd87, 8'd110, 8'd97, 8'd154, 8'd172, 8'd121, 8'd173, 8'd149, 8'd190, 8'd102, 8'd101, 8'd139, 8'd93, 8'd139, 8'd88, 8'd158, 8'd78, 8'd50, 8'd127, 8'd124, 8'd112, 8'd129, 8'd120, 8'd117, 8'd153, 8'd71, 8'd148, 8'd122, 8'd58, 8'd76, 8'd69, 8'd154, 8'd125, 8'd144, 8'd143, 8'd138, 8'd88, 8'd129, 8'd143, 8'd181, 8'd146, 8'd153, 8'd116, 8'd86, 8'd111, 8'd103, 8'd129, 8'd35, 8'd123, 8'd112, 8'd78, 8'd106, 8'd125, 8'd75, 8'd165, 8'd152, 8'd64, 8'd122, 8'd63, 8'd105, 8'd147, 8'd102, 8'd118, 8'd162, 8'd108, 8'd141, 8'd96, 8'd127, 8'd101, 8'd103, 8'd156, 8'd106, 8'd110, 8'd133, 8'd62, 8'd120, 8'd82, 8'd147, 8'd107, 8'd103, 8'd135, 8'd132, 8'd80, 8'd153, 8'd92, 8'd105, 8'd44, 8'd81, 8'd62, 8'd99, 8'd113, 8'd125, 8'd148, 8'd86, 8'd157, 8'd174, 8'd79, 8'd79, 8'd132, 8'd141, 8'd125, 8'd84, 8'd42, 8'd45, 8'd125, 8'd143, 8'd146, 8'd104, 8'd137, 8'd101, 8'd151, 8'd105, 8'd61, 8'd31, 8'd49, 8'd100, 8'd108, 8'd53, 8'd74, 8'd134, 8'd85, 8'd144, 8'd117, 8'd121, 8'd154, 8'd171, 8'd85, 8'd112, 8'd117, 8'd106, 8'd103, 8'd150, 8'd86, 8'd169, 8'd99, 8'd114, 8'd124, 8'd110, 8'd94, 8'd76, 8'd121, 8'd69, 8'd105, 8'd57, 8'd43, 8'd53, 8'd115, 8'd123, 8'd74, 8'd99, 8'd163, 8'd115, 8'd138, 8'd156, 8'd62, 8'd112, 8'd75, 8'd91, 8'd57, 8'd76, 8'd132, 8'd94, 8'd101, 8'd109, 8'd169, 8'd89, 8'd146, 8'd173, 8'd80, 8'd47, 8'd27, 8'd75, 8'd89, 8'd91, 8'd112, 8'd87, 8'd95, 8'd146, 8'd182, 8'd138, 8'd107, 8'd158, 8'd142, 8'd143, 8'd102, 8'd133, 8'd95, 8'd161, 8'd175, 8'd154, 8'd140, 8'd190, 8'd147, 8'd118, 8'd101, 8'd115, 8'd75, 8'd130, 8'd97, 8'd110, 8'd127, 8'd109, 8'd171, 8'd138, 8'd139, 8'd150, 8'd145, 8'd156, 8'd123, 8'd78, 8'd95, 8'd119, 8'd72, 8'd110, 8'd99, 8'd168, 8'd153, 8'd124, 8'd112, 8'd117, 8'd152, 8'd116, 8'd116, 8'd106, 8'd120, 8'd135, 8'd147, 8'd104, 8'd97, 8'd108, 8'd164, 8'd175, 8'd185, 8'd123, 8'd168, 8'd158, 8'd103, 8'd104, 8'd94, 8'd93, 8'd67, 8'd126, 8'd167, 8'd173, 8'd182, 8'd158, 8'd182, 8'd147, 8'd108, 8'd163, 8'd187, 8'd155, 8'd118, 8'd99, 8'd88, 8'd105, 8'd122, 8'd182, 8'd92, 8'd166, 8'd173, 8'd155, 8'd146, 8'd94, 8'd101, 8'd149, 8'd101, 8'd65, 8'd151, 8'd114, 8'd169, 8'd153, 8'd130, 8'd159, 8'd155, 8'd192, 8'd196, 8'd184, 8'd188, 8'd182, 8'd76, 8'd131, 8'd145, 8'd87, 8'd101, 8'd159, 8'd177, 8'd89, 8'd78, 8'd106, 8'd131, 8'd168, 8'd119, 8'd82, 8'd79, 8'd60, 8'd141, 8'd105, 8'd136, 8'd98, 8'd88, 8'd148, 8'd112, 8'd148, 8'd150, 8'd177, 8'd171, 8'd182, 8'd73, 8'd65, 8'd83, 8'd102, 8'd90, 8'd96, 8'd134, 8'd105, 8'd142, 8'd97, 8'd173, 8'd103, 8'd135, 8'd164, 8'd141, 8'd47, 8'd39, 8'd97, 8'd69, 8'd99, 8'd161, 8'd107, 8'd209, 8'd120, 8'd187, 8'd204, 8'd142, 8'd115, 8'd90, 8'd144, 8'd97, 8'd119, 8'd111, 8'd101, 8'd65, 8'd114, 8'd103, 8'd118, 8'd112, 8'd167, 8'd111, 8'd163, 8'd91, 8'd79, 8'd69, 8'd10, 8'd87, 8'd78, 8'd145, 8'd158, 8'd164, 8'd198, 8'd198, 8'd118, 8'd166, 8'd173, 8'd94, 8'd123, 8'd102, 8'd47, 8'd112, 8'd41, 8'd54, 8'd70, 8'd77, 8'd123, 8'd166, 8'd85, 8'd90, 8'd122, 8'd85, 8'd65, 8'd93, 8'd44, 8'd56, 8'd117, 8'd77, 8'd152, 8'd165, 8'd149, 8'd156, 8'd172, 8'd168, 8'd94, 8'd151, 8'd79, 8'd37, 8'd43, 8'd60, 8'd133, 8'd84, 8'd96, 8'd97, 8'd165, 8'd168, 8'd155, 8'd109, 8'd135, 8'd72, 8'd117, 8'd30, 8'd14, 8'd50, 8'd129, 8'd85, 8'd116, 8'd175, 8'd174, 8'd126, 8'd117, 8'd101, 8'd89, 8'd131, 8'd124, 8'd62, 8'd127, 8'd144, 8'd84, 8'd147, 8'd160, 8'd164, 8'd168, 8'd187, 8'd94, 8'd126, 8'd157, 8'd84, 8'd137, 8'd110, 8'd52, 8'd87, 8'd145, 8'd98, 8'd101, 8'd76, 8'd158, 8'd165, 8'd155, 8'd166, 8'd149, 8'd130, 8'd141, 8'd112, 8'd102, 8'd164, 8'd133, 8'd152, 8'd125, 8'd118, 8'd113, 8'd166, 8'd70, 8'd181, 8'd89, 8'd105, 8'd134, 8'd57, 8'd101, 8'd128, 8'd94, 8'd148, 8'd85, 8'd102, 8'd106, 8'd157, 8'd89, 8'd163, 8'd106, 8'd96, 8'd155, 8'd121, 8'd88, 8'd85, 8'd111, 8'd159, 8'd110, 8'd188, 8'd173, 8'd119, 8'd90, 8'd89, 8'd148, 8'd154, 8'd92, 8'd127, 8'd92, 8'd104, 8'd147, 8'd85, 8'd147, 8'd85, 8'd112, 8'd81, 8'd77, 8'd133, 8'd110, 8'd128, 8'd91, 8'd103, 8'd106, 8'd101, 8'd111, 8'd178, 8'd112, 8'd185, 8'd150, 8'd107, 8'd145, 8'd143, 8'd73, 8'd138, 8'd118, 8'd137, 8'd150, 8'd88, 8'd99, 8'd67, 8'd117, 8'd125, 8'd119, 8'd146, 8'd120, 8'd57, 8'd158, 8'd114, 8'd119, 8'd102, 8'd75, 8'd79, 8'd165, 8'd105, 8'd111, 8'd144, 8'd115, 8'd105, 8'd151, 8'd80, 8'd112, 8'd114, 8'd97, 8'd121, 8'd97, 8'd89, 8'd144, 8'd98, 8'd145, 8'd123, 8'd88, 8'd115, 8'd84, 8'd156, 8'd114, 8'd80, 8'd155, 8'd148, 8'd58, 8'd70, 8'd146, 8'd110, 8'd98, 8'd142, 8'd155, 8'd89, 8'd132, 8'd144, 8'd131, 8'd105, 8'd134, 8'd149, 8'd155, 8'd80, 8'd66, 8'd141, 8'd81, 8'd157, 8'd82, 8'd157, 8'd101, 8'd141, 8'd127, 8'd131, 8'd111, 8'd41, 8'd68, 8'd97, 8'd88, 8'd86, 8'd63, 8'd165, 8'd65, 8'd145, 8'd113, 8'd94, 8'd86, 8'd145, 8'd89, 8'd75, 8'd146, 8'd89, 8'd66, 8'd112, 8'd120, 8'd105, 8'd118, 8'd111, 8'd119, 8'd111, 8'd142, 8'd59, 8'd103, 8'd61, 8'd146, 8'd93, 8'd94, 8'd80, 8'd127, 8'd145, 8'd107, 8'd106, 8'd98, 8'd94, 8'd170, 8'd104, 8'd80, 8'd80, 8'd152, 8'd115, 8'd84, 8'd130, 8'd123, 8'd132, 8'd122, 8'd150, 8'd84, 8'd120, 8'd154, 8'd124, 8'd69, 8'd144, 8'd78, 8'd88, 8'd158, 8'd168, 8'd123, 8'd156, 8'd139, 8'd164, 8'd144, 8'd86, 8'd70})
) cell_0_54 (
    .clk(clk),
    .input_index(index_0_53_54),
    .input_value(value_0_53_54),
    .input_result(result_0_53_54),
    .input_enable(enable_0_53_54),
    .output_index(index_0_54_55),
    .output_value(value_0_54_55),
    .output_result(result_0_54_55),
    .output_enable(enable_0_54_55)
);

wire [10-1:0] index_0_55_56;
wire [`DATA_WIDTH-1:0] value_0_55_56;
wire [`DATA_WIDTH*4:0] result_0_55_56;
wire enable_0_55_56;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd155, 8'd80, 8'd140, 8'd99, 8'd94, 8'd109, 8'd123, 8'd149, 8'd191, 8'd126, 8'd168, 8'd164, 8'd164, 8'd140, 8'd204, 8'd135, 8'd185, 8'd117, 8'd88, 8'd133, 8'd161, 8'd158, 8'd136, 8'd85, 8'd94, 8'd164, 8'd101, 8'd145, 8'd145, 8'd76, 8'd87, 8'd102, 8'd80, 8'd149, 8'd114, 8'd92, 8'd149, 8'd172, 8'd178, 8'd122, 8'd105, 8'd107, 8'd112, 8'd121, 8'd132, 8'd86, 8'd91, 8'd102, 8'd111, 8'd77, 8'd100, 8'd147, 8'd71, 8'd128, 8'd160, 8'd131, 8'd114, 8'd160, 8'd150, 8'd94, 8'd159, 8'd132, 8'd89, 8'd118, 8'd151, 8'd154, 8'd101, 8'd103, 8'd143, 8'd133, 8'd137, 8'd138, 8'd204, 8'd120, 8'd144, 8'd132, 8'd135, 8'd121, 8'd136, 8'd111, 8'd122, 8'd91, 8'd87, 8'd87, 8'd76, 8'd148, 8'd94, 8'd155, 8'd118, 8'd164, 8'd130, 8'd136, 8'd160, 8'd151, 8'd170, 8'd155, 8'd76, 8'd83, 8'd83, 8'd133, 8'd82, 8'd126, 8'd173, 8'd95, 8'd178, 8'd110, 8'd200, 8'd114, 8'd141, 8'd80, 8'd157, 8'd92, 8'd137, 8'd86, 8'd91, 8'd114, 8'd119, 8'd106, 8'd110, 8'd88, 8'd117, 8'd120, 8'd150, 8'd134, 8'd146, 8'd103, 8'd110, 8'd78, 8'd148, 8'd76, 8'd82, 8'd117, 8'd126, 8'd132, 8'd124, 8'd164, 8'd186, 8'd164, 8'd134, 8'd92, 8'd106, 8'd122, 8'd127, 8'd96, 8'd142, 8'd168, 8'd109, 8'd92, 8'd119, 8'd107, 8'd76, 8'd162, 8'd151, 8'd97, 8'd79, 8'd142, 8'd156, 8'd128, 8'd124, 8'd92, 8'd141, 8'd152, 8'd111, 8'd122, 8'd124, 8'd96, 8'd140, 8'd118, 8'd68, 8'd156, 8'd138, 8'd124, 8'd143, 8'd150, 8'd119, 8'd98, 8'd108, 8'd98, 8'd106, 8'd97, 8'd90, 8'd182, 8'd153, 8'd93, 8'd173, 8'd161, 8'd148, 8'd162, 8'd190, 8'd153, 8'd132, 8'd161, 8'd143, 8'd178, 8'd78, 8'd148, 8'd174, 8'd176, 8'd152, 8'd137, 8'd146, 8'd142, 8'd103, 8'd123, 8'd127, 8'd124, 8'd142, 8'd133, 8'd188, 8'd152, 8'd188, 8'd171, 8'd119, 8'd129, 8'd149, 8'd144, 8'd157, 8'd98, 8'd158, 8'd193, 8'd210, 8'd100, 8'd96, 8'd128, 8'd135, 8'd179, 8'd128, 8'd146, 8'd178, 8'd135, 8'd152, 8'd122, 8'd182, 8'd133, 8'd175, 8'd184, 8'd185, 8'd191, 8'd173, 8'd169, 8'd135, 8'd104, 8'd177, 8'd124, 8'd174, 8'd115, 8'd126, 8'd196, 8'd147, 8'd99, 8'd99, 8'd98, 8'd163, 8'd121, 8'd158, 8'd178, 8'd141, 8'd186, 8'd152, 8'd146, 8'd125, 8'd178, 8'd147, 8'd89, 8'd72, 8'd161, 8'd142, 8'd135, 8'd120, 8'd88, 8'd84, 8'd47, 8'd89, 8'd97, 8'd119, 8'd136, 8'd181, 8'd147, 8'd177, 8'd125, 8'd155, 8'd183, 8'd158, 8'd173, 8'd158, 8'd111, 8'd158, 8'd137, 8'd145, 8'd155, 8'd78, 8'd124, 8'd116, 8'd102, 8'd89, 8'd99, 8'd92, 8'd56, 8'd44, 8'd109, 8'd120, 8'd123, 8'd159, 8'd211, 8'd141, 8'd171, 8'd135, 8'd81, 8'd168, 8'd160, 8'd187, 8'd185, 8'd140, 8'd139, 8'd124, 8'd103, 8'd115, 8'd89, 8'd96, 8'd97, 8'd64, 8'd159, 8'd140, 8'd131, 8'd124, 8'd133, 8'd107, 8'd68, 8'd89, 8'd118, 8'd105, 8'd114, 8'd136, 8'd174, 8'd82, 8'd154, 8'd177, 8'd170, 8'd173, 8'd131, 8'd161, 8'd90, 8'd136, 8'd73, 8'd146, 8'd124, 8'd110, 8'd90, 8'd84, 8'd128, 8'd110, 8'd134, 8'd108, 8'd55, 8'd65, 8'd82, 8'd111, 8'd48, 8'd126, 8'd130, 8'd94, 8'd137, 8'd106, 8'd89, 8'd142, 8'd140, 8'd103, 8'd99, 8'd108, 8'd130, 8'd111, 8'd141, 8'd124, 8'd108, 8'd130, 8'd72, 8'd125, 8'd157, 8'd113, 8'd155, 8'd100, 8'd112, 8'd69, 8'd69, 8'd56, 8'd61, 8'd98, 8'd99, 8'd100, 8'd145, 8'd154, 8'd176, 8'd85, 8'd194, 8'd130, 8'd122, 8'd31, 8'd16, 8'd76, 8'd35, 8'd104, 8'd134, 8'd70, 8'd97, 8'd185, 8'd130, 8'd153, 8'd127, 8'd74, 8'd61, 8'd65, 8'd30, 8'd95, 8'd62, 8'd126, 8'd154, 8'd152, 8'd117, 8'd144, 8'd106, 8'd172, 8'd98, 8'd145, 8'd50, 8'd100, 8'd7, 8'd55, 8'd72, 8'd47, 8'd86, 8'd126, 8'd107, 8'd97, 8'd117, 8'd92, 8'd107, 8'd57, 8'd40, 8'd34, 8'd99, 8'd15, 8'd110, 8'd139, 8'd111, 8'd123, 8'd151, 8'd126, 8'd104, 8'd140, 8'd112, 8'd152, 8'd93, 8'd46, 8'd87, 8'd33, 8'd54, 8'd145, 8'd132, 8'd94, 8'd105, 8'd188, 8'd203, 8'd114, 8'd31, 8'd38, 8'd111, 8'd65, 8'd93, 8'd115, 8'd51, 8'd121, 8'd114, 8'd122, 8'd198, 8'd115, 8'd135, 8'd137, 8'd204, 8'd143, 8'd130, 8'd51, 8'd102, 8'd81, 8'd85, 8'd93, 8'd55, 8'd152, 8'd101, 8'd213, 8'd194, 8'd147, 8'd50, 8'd112, 8'd70, 8'd90, 8'd98, 8'd95, 8'd168, 8'd161, 8'd112, 8'd148, 8'd197, 8'd134, 8'd103, 8'd123, 8'd145, 8'd193, 8'd72, 8'd113, 8'd38, 8'd129, 8'd63, 8'd112, 8'd127, 8'd66, 8'd152, 8'd218, 8'd147, 8'd150, 8'd116, 8'd83, 8'd139, 8'd104, 8'd112, 8'd99, 8'd149, 8'd166, 8'd170, 8'd154, 8'd166, 8'd115, 8'd121, 8'd88, 8'd134, 8'd133, 8'd56, 8'd8, 8'd93, 8'd92, 8'd69, 8'd133, 8'd91, 8'd106, 8'd108, 8'd154, 8'd177, 8'd160, 8'd182, 8'd128, 8'd111, 8'd124, 8'd98, 8'd178, 8'd114, 8'd151, 8'd123, 8'd138, 8'd133, 8'd133, 8'd82, 8'd100, 8'd116, 8'd159, 8'd24, 8'd49, 8'd38, 8'd124, 8'd111, 8'd151, 8'd65, 8'd131, 8'd197, 8'd156, 8'd221, 8'd123, 8'd153, 8'd160, 8'd170, 8'd120, 8'd125, 8'd165, 8'd137, 8'd132, 8'd172, 8'd101, 8'd176, 8'd144, 8'd137, 8'd101, 8'd81, 8'd87, 8'd103, 8'd44, 8'd51, 8'd113, 8'd56, 8'd122, 8'd138, 8'd120, 8'd185, 8'd176, 8'd181, 8'd112, 8'd132, 8'd138, 8'd93, 8'd117, 8'd85, 8'd95, 8'd165, 8'd148, 8'd146, 8'd126, 8'd167, 8'd86, 8'd128, 8'd151, 8'd101, 8'd69, 8'd61, 8'd41, 8'd88, 8'd149, 8'd62, 8'd119, 8'd152, 8'd103, 8'd81, 8'd114, 8'd97, 8'd97, 8'd108, 8'd106, 8'd109, 8'd87, 8'd148, 8'd146, 8'd138, 8'd104, 8'd108, 8'd177, 8'd136, 8'd110, 8'd76, 8'd119, 8'd166, 8'd165, 8'd107, 8'd104, 8'd87, 8'd103, 8'd118, 8'd96, 8'd172, 8'd177, 8'd165, 8'd159, 8'd119, 8'd171, 8'd148, 8'd198, 8'd207, 8'd140, 8'd189, 8'd195, 8'd117, 8'd100, 8'd170, 8'd160, 8'd90, 8'd127, 8'd148, 8'd94, 8'd94, 8'd127, 8'd84, 8'd143, 8'd127, 8'd112, 8'd155, 8'd152, 8'd216, 8'd154, 8'd213, 8'd196, 8'd203, 8'd255, 8'd183, 8'd164, 8'd194, 8'd214, 8'd207, 8'd162, 8'd165, 8'd85, 8'd121, 8'd100, 8'd142, 8'd107, 8'd119, 8'd133, 8'd145, 8'd140, 8'd179, 8'd152, 8'd105, 8'd178, 8'd137, 8'd132, 8'd160, 8'd187, 8'd237, 8'd247, 8'd207, 8'd210, 8'd210, 8'd191, 8'd129, 8'd169, 8'd183, 8'd137, 8'd161, 8'd157, 8'd140, 8'd97, 8'd144, 8'd86, 8'd126, 8'd70, 8'd102, 8'd118, 8'd116, 8'd112, 8'd108, 8'd134, 8'd132, 8'd108, 8'd113, 8'd118, 8'd136, 8'd127, 8'd122, 8'd158, 8'd159, 8'd154, 8'd183, 8'd122, 8'd180, 8'd121, 8'd114, 8'd90, 8'd75, 8'd79, 8'd160, 8'd162, 8'd104, 8'd137, 8'd167, 8'd156, 8'd128, 8'd117, 8'd108, 8'd150, 8'd166, 8'd168, 8'd105, 8'd162, 8'd144, 8'd141, 8'd103, 8'd148, 8'd119, 8'd78, 8'd77, 8'd137, 8'd125, 8'd146, 8'd98, 8'd120, 8'd117, 8'd140, 8'd132, 8'd122, 8'd107})
) cell_0_55 (
    .clk(clk),
    .input_index(index_0_54_55),
    .input_value(value_0_54_55),
    .input_result(result_0_54_55),
    .input_enable(enable_0_54_55),
    .output_index(index_0_55_56),
    .output_value(value_0_55_56),
    .output_result(result_0_55_56),
    .output_enable(enable_0_55_56)
);

wire [10-1:0] index_0_56_57;
wire [`DATA_WIDTH-1:0] value_0_56_57;
wire [`DATA_WIDTH*4:0] result_0_56_57;
wire enable_0_56_57;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd151, 8'd109, 8'd107, 8'd91, 8'd96, 8'd122, 8'd86, 8'd107, 8'd125, 8'd100, 8'd126, 8'd62, 8'd85, 8'd74, 8'd43, 8'd70, 8'd156, 8'd100, 8'd94, 8'd146, 8'd76, 8'd99, 8'd126, 8'd90, 8'd138, 8'd104, 8'd80, 8'd109, 8'd102, 8'd80, 8'd96, 8'd150, 8'd91, 8'd129, 8'd110, 8'd94, 8'd103, 8'd53, 8'd144, 8'd111, 8'd128, 8'd103, 8'd61, 8'd57, 8'd126, 8'd102, 8'd78, 8'd96, 8'd87, 8'd159, 8'd146, 8'd116, 8'd130, 8'd100, 8'd111, 8'd122, 8'd82, 8'd127, 8'd69, 8'd162, 8'd129, 8'd131, 8'd130, 8'd156, 8'd135, 8'd147, 8'd116, 8'd142, 8'd61, 8'd74, 8'd52, 8'd143, 8'd120, 8'd100, 8'd76, 8'd73, 8'd119, 8'd120, 8'd143, 8'd72, 8'd58, 8'd95, 8'd148, 8'd114, 8'd96, 8'd77, 8'd154, 8'd165, 8'd94, 8'd139, 8'd184, 8'd141, 8'd179, 8'd164, 8'd122, 8'd166, 8'd125, 8'd156, 8'd156, 8'd143, 8'd76, 8'd102, 8'd82, 8'd73, 8'd92, 8'd85, 8'd53, 8'd87, 8'd59, 8'd77, 8'd109, 8'd108, 8'd169, 8'd86, 8'd127, 8'd151, 8'd101, 8'd117, 8'd172, 8'd136, 8'd152, 8'd161, 8'd126, 8'd167, 8'd102, 8'd97, 8'd156, 8'd167, 8'd126, 8'd71, 8'd111, 8'd157, 8'd80, 8'd100, 8'd127, 8'd95, 8'd72, 8'd114, 8'd142, 8'd83, 8'd115, 8'd146, 8'd96, 8'd93, 8'd101, 8'd135, 8'd121, 8'd98, 8'd99, 8'd170, 8'd108, 8'd166, 8'd133, 8'd140, 8'd87, 8'd107, 8'd80, 8'd146, 8'd143, 8'd75, 8'd75, 8'd63, 8'd57, 8'd138, 8'd136, 8'd119, 8'd137, 8'd151, 8'd149, 8'd96, 8'd98, 8'd84, 8'd119, 8'd145, 8'd192, 8'd112, 8'd170, 8'd129, 8'd103, 8'd149, 8'd154, 8'd129, 8'd109, 8'd88, 8'd100, 8'd113, 8'd134, 8'd111, 8'd73, 8'd101, 8'd74, 8'd140, 8'd137, 8'd102, 8'd147, 8'd94, 8'd126, 8'd98, 8'd67, 8'd112, 8'd123, 8'd164, 8'd141, 8'd134, 8'd160, 8'd128, 8'd123, 8'd126, 8'd122, 8'd137, 8'd74, 8'd133, 8'd77, 8'd50, 8'd116, 8'd137, 8'd170, 8'd162, 8'd132, 8'd93, 8'd63, 8'd113, 8'd99, 8'd125, 8'd87, 8'd110, 8'd70, 8'd74, 8'd170, 8'd125, 8'd152, 8'd84, 8'd164, 8'd177, 8'd158, 8'd106, 8'd154, 8'd96, 8'd74, 8'd110, 8'd125, 8'd147, 8'd75, 8'd103, 8'd137, 8'd104, 8'd93, 8'd111, 8'd118, 8'd132, 8'd145, 8'd148, 8'd122, 8'd114, 8'd15, 8'd112, 8'd155, 8'd141, 8'd105, 8'd72, 8'd157, 8'd138, 8'd161, 8'd130, 8'd87, 8'd132, 8'd56, 8'd72, 8'd174, 8'd173, 8'd128, 8'd186, 8'd157, 8'd71, 8'd54, 8'd67, 8'd82, 8'd99, 8'd127, 8'd70, 8'd135, 8'd89, 8'd107, 8'd61, 8'd69, 8'd122, 8'd70, 8'd132, 8'd70, 8'd81, 8'd162, 8'd111, 8'd163, 8'd139, 8'd129, 8'd135, 8'd193, 8'd112, 8'd113, 8'd117, 8'd189, 8'd70, 8'd112, 8'd115, 8'd107, 8'd156, 8'd88, 8'd102, 8'd134, 8'd83, 8'd130, 8'd125, 8'd48, 8'd64, 8'd144, 8'd141, 8'd62, 8'd82, 8'd82, 8'd136, 8'd180, 8'd115, 8'd128, 8'd113, 8'd136, 8'd177, 8'd122, 8'd124, 8'd87, 8'd96, 8'd80, 8'd92, 8'd118, 8'd79, 8'd157, 8'd141, 8'd78, 8'd141, 8'd129, 8'd72, 8'd90, 8'd113, 8'd125, 8'd75, 8'd138, 8'd152, 8'd127, 8'd167, 8'd116, 8'd121, 8'd173, 8'd144, 8'd206, 8'd164, 8'd194, 8'd119, 8'd142, 8'd142, 8'd84, 8'd127, 8'd114, 8'd144, 8'd159, 8'd76, 8'd109, 8'd93, 8'd75, 8'd51, 8'd68, 8'd87, 8'd143, 8'd147, 8'd104, 8'd124, 8'd124, 8'd190, 8'd144, 8'd119, 8'd167, 8'd230, 8'd228, 8'd149, 8'd186, 8'd134, 8'd88, 8'd165, 8'd116, 8'd136, 8'd63, 8'd66, 8'd107, 8'd90, 8'd159, 8'd149, 8'd132, 8'd92, 8'd141, 8'd99, 8'd152, 8'd163, 8'd158, 8'd82, 8'd151, 8'd96, 8'd143, 8'd167, 8'd239, 8'd221, 8'd213, 8'd193, 8'd114, 8'd157, 8'd172, 8'd133, 8'd171, 8'd84, 8'd101, 8'd99, 8'd132, 8'd114, 8'd75, 8'd66, 8'd94, 8'd144, 8'd190, 8'd183, 8'd125, 8'd117, 8'd118, 8'd97, 8'd141, 8'd81, 8'd158, 8'd158, 8'd150, 8'd158, 8'd213, 8'd157, 8'd154, 8'd181, 8'd125, 8'd111, 8'd157, 8'd78, 8'd71, 8'd118, 8'd149, 8'd132, 8'd135, 8'd123, 8'd118, 8'd140, 8'd120, 8'd176, 8'd95, 8'd161, 8'd84, 8'd128, 8'd117, 8'd62, 8'd90, 8'd98, 8'd169, 8'd158, 8'd190, 8'd171, 8'd184, 8'd170, 8'd174, 8'd112, 8'd131, 8'd91, 8'd66, 8'd54, 8'd71, 8'd94, 8'd123, 8'd142, 8'd136, 8'd80, 8'd82, 8'd102, 8'd123, 8'd111, 8'd83, 8'd100, 8'd69, 8'd97, 8'd74, 8'd101, 8'd86, 8'd167, 8'd131, 8'd137, 8'd165, 8'd148, 8'd106, 8'd126, 8'd142, 8'd56, 8'd102, 8'd45, 8'd80, 8'd69, 8'd74, 8'd98, 8'd126, 8'd141, 8'd165, 8'd108, 8'd125, 8'd145, 8'd92, 8'd148, 8'd65, 8'd90, 8'd52, 8'd58, 8'd55, 8'd115, 8'd115, 8'd123, 8'd90, 8'd103, 8'd163, 8'd114, 8'd123, 8'd123, 8'd91, 8'd72, 8'd122, 8'd101, 8'd131, 8'd172, 8'd174, 8'd127, 8'd157, 8'd153, 8'd138, 8'd126, 8'd109, 8'd96, 8'd84, 8'd88, 8'd125, 8'd107, 8'd56, 8'd58, 8'd109, 8'd143, 8'd84, 8'd67, 8'd138, 8'd150, 8'd70, 8'd69, 8'd89, 8'd64, 8'd72, 8'd124, 8'd116, 8'd151, 8'd150, 8'd199, 8'd152, 8'd127, 8'd146, 8'd137, 8'd102, 8'd76, 8'd103, 8'd153, 8'd82, 8'd76, 8'd89, 8'd133, 8'd66, 8'd116, 8'd136, 8'd91, 8'd61, 8'd129, 8'd83, 8'd98, 8'd50, 8'd76, 8'd102, 8'd74, 8'd132, 8'd152, 8'd127, 8'd147, 8'd180, 8'd140, 8'd150, 8'd107, 8'd166, 8'd111, 8'd150, 8'd141, 8'd88, 8'd128, 8'd106, 8'd85, 8'd142, 8'd103, 8'd119, 8'd114, 8'd105, 8'd65, 8'd101, 8'd130, 8'd57, 8'd139, 8'd65, 8'd132, 8'd167, 8'd94, 8'd138, 8'd81, 8'd97, 8'd160, 8'd132, 8'd111, 8'd174, 8'd178, 8'd114, 8'd93, 8'd180, 8'd143, 8'd151, 8'd121, 8'd138, 8'd150, 8'd161, 8'd78, 8'd73, 8'd101, 8'd153, 8'd89, 8'd153, 8'd80, 8'd79, 8'd74, 8'd103, 8'd168, 8'd149, 8'd124, 8'd72, 8'd86, 8'd90, 8'd114, 8'd122, 8'd60, 8'd138, 8'd138, 8'd95, 8'd85, 8'd97, 8'd72, 8'd75, 8'd86, 8'd86, 8'd108, 8'd150, 8'd129, 8'd171, 8'd86, 8'd120, 8'd109, 8'd123, 8'd125, 8'd148, 8'd128, 8'd137, 8'd92, 8'd131, 8'd125, 8'd142, 8'd65, 8'd108, 8'd50, 8'd57, 8'd75, 8'd101, 8'd65, 8'd18, 8'd73, 8'd113, 8'd120, 8'd90, 8'd110, 8'd84, 8'd98, 8'd99, 8'd92, 8'd97, 8'd124, 8'd152, 8'd86, 8'd109, 8'd73, 8'd95, 8'd115, 8'd67, 8'd133, 8'd98, 8'd69, 8'd105, 8'd146, 8'd42, 8'd123, 8'd75, 8'd120, 8'd74, 8'd88, 8'd95, 8'd53, 8'd105, 8'd68, 8'd123, 8'd112, 8'd141, 8'd146, 8'd102, 8'd99, 8'd150, 8'd155, 8'd142, 8'd118, 8'd139, 8'd79, 8'd104, 8'd126, 8'd118, 8'd60, 8'd90, 8'd64, 8'd132, 8'd125, 8'd54, 8'd106, 8'd64, 8'd67, 8'd98, 8'd78, 8'd127, 8'd129, 8'd112, 8'd155, 8'd128, 8'd164, 8'd88, 8'd115, 8'd121, 8'd88, 8'd119, 8'd80, 8'd79, 8'd75, 8'd85, 8'd78, 8'd161, 8'd137, 8'd127, 8'd114, 8'd110, 8'd70, 8'd129, 8'd166, 8'd100, 8'd70, 8'd114, 8'd141, 8'd120, 8'd78, 8'd82, 8'd136, 8'd167, 8'd114, 8'd106, 8'd116, 8'd108, 8'd118})
) cell_0_56 (
    .clk(clk),
    .input_index(index_0_55_56),
    .input_value(value_0_55_56),
    .input_result(result_0_55_56),
    .input_enable(enable_0_55_56),
    .output_index(index_0_56_57),
    .output_value(value_0_56_57),
    .output_result(result_0_56_57),
    .output_enable(enable_0_56_57)
);

wire [10-1:0] index_0_57_58;
wire [`DATA_WIDTH-1:0] value_0_57_58;
wire [`DATA_WIDTH*4:0] result_0_57_58;
wire enable_0_57_58;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd101, 8'd123, 8'd124, 8'd78, 8'd72, 8'd103, 8'd158, 8'd164, 8'd78, 8'd68, 8'd70, 8'd148, 8'd148, 8'd85, 8'd83, 8'd134, 8'd148, 8'd63, 8'd142, 8'd75, 8'd153, 8'd125, 8'd77, 8'd120, 8'd128, 8'd152, 8'd114, 8'd151, 8'd152, 8'd121, 8'd155, 8'd115, 8'd153, 8'd135, 8'd85, 8'd131, 8'd154, 8'd84, 8'd73, 8'd90, 8'd61, 8'd157, 8'd155, 8'd142, 8'd134, 8'd102, 8'd89, 8'd134, 8'd119, 8'd87, 8'd76, 8'd130, 8'd103, 8'd88, 8'd125, 8'd146, 8'd127, 8'd150, 8'd120, 8'd79, 8'd95, 8'd122, 8'd164, 8'd173, 8'd81, 8'd125, 8'd104, 8'd92, 8'd75, 8'd118, 8'd79, 8'd143, 8'd125, 8'd126, 8'd61, 8'd81, 8'd54, 8'd137, 8'd85, 8'd108, 8'd57, 8'd92, 8'd118, 8'd120, 8'd170, 8'd107, 8'd92, 8'd71, 8'd159, 8'd132, 8'd168, 8'd94, 8'd122, 8'd174, 8'd156, 8'd111, 8'd177, 8'd133, 8'd82, 8'd127, 8'd100, 8'd89, 8'd108, 8'd154, 8'd127, 8'd32, 8'd91, 8'd73, 8'd90, 8'd99, 8'd149, 8'd85, 8'd155, 8'd79, 8'd102, 8'd150, 8'd79, 8'd136, 8'd170, 8'd107, 8'd144, 8'd89, 8'd109, 8'd99, 8'd126, 8'd92, 8'd91, 8'd123, 8'd168, 8'd113, 8'd136, 8'd103, 8'd157, 8'd110, 8'd55, 8'd108, 8'd71, 8'd85, 8'd133, 8'd145, 8'd119, 8'd134, 8'd65, 8'd88, 8'd113, 8'd145, 8'd138, 8'd149, 8'd164, 8'd92, 8'd166, 8'd76, 8'd133, 8'd91, 8'd157, 8'd143, 8'd88, 8'd117, 8'd66, 8'd158, 8'd140, 8'd79, 8'd114, 8'd100, 8'd142, 8'd86, 8'd135, 8'd140, 8'd143, 8'd119, 8'd64, 8'd87, 8'd143, 8'd163, 8'd77, 8'd167, 8'd160, 8'd151, 8'd125, 8'd147, 8'd139, 8'd138, 8'd137, 8'd105, 8'd101, 8'd77, 8'd81, 8'd108, 8'd82, 8'd113, 8'd95, 8'd125, 8'd46, 8'd72, 8'd115, 8'd161, 8'd148, 8'd61, 8'd147, 8'd153, 8'd166, 8'd98, 8'd144, 8'd121, 8'd104, 8'd164, 8'd82, 8'd102, 8'd164, 8'd137, 8'd115, 8'd134, 8'd148, 8'd142, 8'd154, 8'd97, 8'd91, 8'd160, 8'd91, 8'd109, 8'd117, 8'd106, 8'd109, 8'd111, 8'd83, 8'd55, 8'd144, 8'd97, 8'd77, 8'd138, 8'd104, 8'd159, 8'd99, 8'd77, 8'd94, 8'd78, 8'd123, 8'd122, 8'd112, 8'd158, 8'd172, 8'd140, 8'd150, 8'd80, 8'd83, 8'd121, 8'd85, 8'd133, 8'd32, 8'd87, 8'd146, 8'd138, 8'd131, 8'd131, 8'd118, 8'd155, 8'd151, 8'd71, 8'd139, 8'd71, 8'd85, 8'd105, 8'd136, 8'd143, 8'd81, 8'd99, 8'd133, 8'd164, 8'd154, 8'd137, 8'd174, 8'd116, 8'd111, 8'd81, 8'd58, 8'd64, 8'd90, 8'd119, 8'd76, 8'd164, 8'd135, 8'd93, 8'd148, 8'd65, 8'd107, 8'd139, 8'd159, 8'd107, 8'd78, 8'd123, 8'd91, 8'd93, 8'd109, 8'd90, 8'd126, 8'd113, 8'd152, 8'd166, 8'd169, 8'd186, 8'd183, 8'd100, 8'd126, 8'd93, 8'd67, 8'd117, 8'd93, 8'd149, 8'd149, 8'd148, 8'd121, 8'd109, 8'd156, 8'd59, 8'd64, 8'd126, 8'd48, 8'd145, 8'd75, 8'd98, 8'd103, 8'd178, 8'd116, 8'd124, 8'd124, 8'd177, 8'd115, 8'd125, 8'd135, 8'd145, 8'd86, 8'd65, 8'd76, 8'd71, 8'd153, 8'd110, 8'd133, 8'd66, 8'd130, 8'd106, 8'd132, 8'd118, 8'd117, 8'd135, 8'd125, 8'd73, 8'd112, 8'd161, 8'd148, 8'd171, 8'd109, 8'd166, 8'd144, 8'd162, 8'd88, 8'd86, 8'd86, 8'd150, 8'd148, 8'd78, 8'd120, 8'd87, 8'd131, 8'd133, 8'd161, 8'd136, 8'd150, 8'd149, 8'd163, 8'd92, 8'd162, 8'd101, 8'd142, 8'd103, 8'd84, 8'd95, 8'd113, 8'd104, 8'd142, 8'd123, 8'd121, 8'd77, 8'd65, 8'd76, 8'd158, 8'd111, 8'd138, 8'd138, 8'd131, 8'd107, 8'd91, 8'd156, 8'd164, 8'd129, 8'd166, 8'd119, 8'd172, 8'd144, 8'd96, 8'd82, 8'd110, 8'd109, 8'd91, 8'd99, 8'd152, 8'd135, 8'd164, 8'd142, 8'd167, 8'd156, 8'd73, 8'd87, 8'd161, 8'd107, 8'd158, 8'd147, 8'd111, 8'd51, 8'd116, 8'd160, 8'd75, 8'd126, 8'd154, 8'd156, 8'd168, 8'd150, 8'd162, 8'd195, 8'd110, 8'd102, 8'd86, 8'd164, 8'd146, 8'd166, 8'd96, 8'd178, 8'd102, 8'd113, 8'd181, 8'd87, 8'd89, 8'd167, 8'd106, 8'd123, 8'd116, 8'd44, 8'd113, 8'd158, 8'd158, 8'd146, 8'd77, 8'd94, 8'd153, 8'd128, 8'd188, 8'd142, 8'd86, 8'd159, 8'd76, 8'd82, 8'd117, 8'd91, 8'd153, 8'd132, 8'd128, 8'd168, 8'd92, 8'd123, 8'd124, 8'd133, 8'd134, 8'd68, 8'd126, 8'd71, 8'd130, 8'd117, 8'd165, 8'd76, 8'd114, 8'd99, 8'd121, 8'd149, 8'd91, 8'd90, 8'd137, 8'd146, 8'd100, 8'd67, 8'd88, 8'd82, 8'd118, 8'd88, 8'd114, 8'd158, 8'd127, 8'd171, 8'd95, 8'd142, 8'd80, 8'd149, 8'd49, 8'd59, 8'd145, 8'd148, 8'd119, 8'd76, 8'd59, 8'd80, 8'd107, 8'd170, 8'd163, 8'd88, 8'd158, 8'd161, 8'd104, 8'd107, 8'd110, 8'd90, 8'd130, 8'd110, 8'd144, 8'd94, 8'd89, 8'd168, 8'd104, 8'd176, 8'd103, 8'd90, 8'd77, 8'd123, 8'd66, 8'd138, 8'd133, 8'd69, 8'd146, 8'd102, 8'd141, 8'd135, 8'd108, 8'd137, 8'd141, 8'd139, 8'd116, 8'd132, 8'd94, 8'd72, 8'd138, 8'd136, 8'd111, 8'd132, 8'd140, 8'd118, 8'd139, 8'd106, 8'd85, 8'd163, 8'd71, 8'd51, 8'd94, 8'd125, 8'd100, 8'd105, 8'd137, 8'd75, 8'd108, 8'd167, 8'd142, 8'd90, 8'd99, 8'd100, 8'd64, 8'd107, 8'd96, 8'd58, 8'd129, 8'd127, 8'd127, 8'd156, 8'd85, 8'd102, 8'd98, 8'd98, 8'd119, 8'd98, 8'd47, 8'd129, 8'd97, 8'd111, 8'd76, 8'd134, 8'd111, 8'd141, 8'd139, 8'd71, 8'd176, 8'd148, 8'd128, 8'd115, 8'd122, 8'd119, 8'd146, 8'd101, 8'd99, 8'd137, 8'd132, 8'd164, 8'd90, 8'd149, 8'd145, 8'd58, 8'd128, 8'd75, 8'd138, 8'd96, 8'd108, 8'd131, 8'd138, 8'd104, 8'd89, 8'd102, 8'd107, 8'd81, 8'd143, 8'd103, 8'd109, 8'd172, 8'd138, 8'd173, 8'd126, 8'd140, 8'd181, 8'd150, 8'd131, 8'd69, 8'd102, 8'd105, 8'd109, 8'd108, 8'd89, 8'd112, 8'd85, 8'd133, 8'd118, 8'd162, 8'd75, 8'd75, 8'd120, 8'd107, 8'd88, 8'd79, 8'd134, 8'd84, 8'd99, 8'd80, 8'd131, 8'd101, 8'd90, 8'd94, 8'd136, 8'd90, 8'd122, 8'd166, 8'd138, 8'd141, 8'd159, 8'd93, 8'd164, 8'd151, 8'd99, 8'd121, 8'd144, 8'd149, 8'd90, 8'd132, 8'd109, 8'd171, 8'd104, 8'd93, 8'd161, 8'd72, 8'd109, 8'd106, 8'd59, 8'd159, 8'd123, 8'd88, 8'd90, 8'd109, 8'd165, 8'd123, 8'd182, 8'd179, 8'd142, 8'd172, 8'd145, 8'd94, 8'd136, 8'd117, 8'd144, 8'd119, 8'd110, 8'd123, 8'd68, 8'd96, 8'd156, 8'd119, 8'd155, 8'd126, 8'd145, 8'd164, 8'd178, 8'd186, 8'd127, 8'd185, 8'd189, 8'd200, 8'd182, 8'd176, 8'd122, 8'd130, 8'd164, 8'd91, 8'd119, 8'd124, 8'd103, 8'd87, 8'd94, 8'd126, 8'd112, 8'd132, 8'd149, 8'd124, 8'd121, 8'd106, 8'd145, 8'd135, 8'd122, 8'd141, 8'd148, 8'd92, 8'd161, 8'd91, 8'd188, 8'd187, 8'd171, 8'd183, 8'd129, 8'd91, 8'd99, 8'd104, 8'd167, 8'd131, 8'd143, 8'd84, 8'd159, 8'd123, 8'd76, 8'd85, 8'd87, 8'd155, 8'd158, 8'd86, 8'd118, 8'd90, 8'd158, 8'd128, 8'd96, 8'd137, 8'd142, 8'd73, 8'd119, 8'd134, 8'd91, 8'd77, 8'd109, 8'd107, 8'd96, 8'd125, 8'd90, 8'd93, 8'd95, 8'd75, 8'd72, 8'd164})
) cell_0_57 (
    .clk(clk),
    .input_index(index_0_56_57),
    .input_value(value_0_56_57),
    .input_result(result_0_56_57),
    .input_enable(enable_0_56_57),
    .output_index(index_0_57_58),
    .output_value(value_0_57_58),
    .output_result(result_0_57_58),
    .output_enable(enable_0_57_58)
);

wire [10-1:0] index_0_58_59;
wire [`DATA_WIDTH-1:0] value_0_58_59;
wire [`DATA_WIDTH*4:0] result_0_58_59;
wire enable_0_58_59;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd147, 8'd154, 8'd118, 8'd141, 8'd102, 8'd91, 8'd106, 8'd117, 8'd150, 8'd104, 8'd112, 8'd144, 8'd75, 8'd114, 8'd134, 8'd124, 8'd77, 8'd67, 8'd136, 8'd87, 8'd104, 8'd151, 8'd79, 8'd94, 8'd120, 8'd118, 8'd111, 8'd127, 8'd134, 8'd109, 8'd70, 8'd88, 8'd77, 8'd109, 8'd157, 8'd165, 8'd173, 8'd130, 8'd101, 8'd75, 8'd116, 8'd93, 8'd145, 8'd93, 8'd126, 8'd146, 8'd88, 8'd132, 8'd126, 8'd128, 8'd123, 8'd181, 8'd79, 8'd76, 8'd163, 8'd104, 8'd73, 8'd105, 8'd154, 8'd81, 8'd104, 8'd135, 8'd95, 8'd183, 8'd113, 8'd144, 8'd92, 8'd102, 8'd157, 8'd138, 8'd117, 8'd161, 8'd91, 8'd166, 8'd182, 8'd126, 8'd181, 8'd107, 8'd145, 8'd161, 8'd122, 8'd144, 8'd162, 8'd85, 8'd126, 8'd85, 8'd64, 8'd138, 8'd91, 8'd134, 8'd172, 8'd87, 8'd114, 8'd75, 8'd142, 8'd108, 8'd80, 8'd130, 8'd59, 8'd153, 8'd127, 8'd126, 8'd133, 8'd95, 8'd119, 8'd176, 8'd152, 8'd116, 8'd129, 8'd124, 8'd113, 8'd163, 8'd85, 8'd116, 8'd68, 8'd64, 8'd117, 8'd75, 8'd92, 8'd165, 8'd120, 8'd111, 8'd117, 8'd136, 8'd136, 8'd138, 8'd137, 8'd165, 8'd157, 8'd106, 8'd131, 8'd143, 8'd172, 8'd92, 8'd126, 8'd144, 8'd75, 8'd166, 8'd119, 8'd118, 8'd111, 8'd145, 8'd125, 8'd90, 8'd80, 8'd124, 8'd91, 8'd70, 8'd108, 8'd65, 8'd133, 8'd63, 8'd144, 8'd136, 8'd106, 8'd115, 8'd141, 8'd112, 8'd129, 8'd95, 8'd108, 8'd168, 8'd139, 8'd87, 8'd93, 8'd143, 8'd146, 8'd150, 8'd132, 8'd141, 8'd97, 8'd150, 8'd93, 8'd146, 8'd81, 8'd103, 8'd78, 8'd123, 8'd108, 8'd95, 8'd97, 8'd142, 8'd77, 8'd77, 8'd71, 8'd113, 8'd121, 8'd135, 8'd134, 8'd147, 8'd144, 8'd146, 8'd90, 8'd152, 8'd158, 8'd106, 8'd133, 8'd139, 8'd96, 8'd103, 8'd94, 8'd117, 8'd144, 8'd81, 8'd137, 8'd139, 8'd67, 8'd96, 8'd66, 8'd103, 8'd102, 8'd59, 8'd81, 8'd107, 8'd40, 8'd55, 8'd99, 8'd83, 8'd150, 8'd71, 8'd70, 8'd128, 8'd102, 8'd166, 8'd132, 8'd129, 8'd80, 8'd95, 8'd73, 8'd123, 8'd84, 8'd116, 8'd117, 8'd92, 8'd83, 8'd123, 8'd60, 8'd61, 8'd99, 8'd88, 8'd67, 8'd81, 8'd125, 8'd64, 8'd103, 8'd75, 8'd100, 8'd104, 8'd61, 8'd107, 8'd78, 8'd119, 8'd145, 8'd142, 8'd45, 8'd75, 8'd113, 8'd144, 8'd120, 8'd143, 8'd65, 8'd121, 8'd141, 8'd87, 8'd79, 8'd65, 8'd68, 8'd75, 8'd44, 8'd129, 8'd155, 8'd166, 8'd92, 8'd67, 8'd79, 8'd94, 8'd68, 8'd75, 8'd146, 8'd160, 8'd136, 8'd49, 8'd29, 8'd64, 8'd64, 8'd85, 8'd65, 8'd121, 8'd106, 8'd109, 8'd165, 8'd149, 8'd136, 8'd127, 8'd66, 8'd119, 8'd78, 8'd143, 8'd139, 8'd107, 8'd169, 8'd136, 8'd97, 8'd77, 8'd104, 8'd141, 8'd171, 8'd77, 8'd109, 8'd78, 8'd104, 8'd54, 8'd132, 8'd104, 8'd80, 8'd103, 8'd119, 8'd173, 8'd93, 8'd158, 8'd103, 8'd85, 8'd113, 8'd77, 8'd85, 8'd169, 8'd119, 8'd118, 8'd130, 8'd125, 8'd127, 8'd103, 8'd93, 8'd88, 8'd147, 8'd159, 8'd125, 8'd93, 8'd131, 8'd135, 8'd94, 8'd172, 8'd127, 8'd103, 8'd158, 8'd97, 8'd96, 8'd133, 8'd169, 8'd133, 8'd134, 8'd134, 8'd117, 8'd92, 8'd172, 8'd143, 8'd129, 8'd127, 8'd131, 8'd153, 8'd77, 8'd143, 8'd141, 8'd83, 8'd126, 8'd123, 8'd51, 8'd66, 8'd147, 8'd102, 8'd94, 8'd110, 8'd121, 8'd145, 8'd149, 8'd152, 8'd109, 8'd132, 8'd116, 8'd112, 8'd88, 8'd151, 8'd162, 8'd103, 8'd154, 8'd181, 8'd194, 8'd177, 8'd98, 8'd61, 8'd121, 8'd97, 8'd100, 8'd32, 8'd78, 8'd87, 8'd126, 8'd150, 8'd158, 8'd116, 8'd147, 8'd167, 8'd132, 8'd109, 8'd116, 8'd176, 8'd98, 8'd165, 8'd128, 8'd141, 8'd185, 8'd108, 8'd155, 8'd141, 8'd122, 8'd136, 8'd136, 8'd60, 8'd82, 8'd87, 8'd84, 8'd120, 8'd59, 8'd178, 8'd202, 8'd185, 8'd144, 8'd121, 8'd147, 8'd100, 8'd142, 8'd116, 8'd153, 8'd134, 8'd85, 8'd161, 8'd176, 8'd139, 8'd146, 8'd160, 8'd186, 8'd152, 8'd179, 8'd92, 8'd77, 8'd60, 8'd55, 8'd130, 8'd67, 8'd126, 8'd49, 8'd68, 8'd105, 8'd148, 8'd105, 8'd162, 8'd185, 8'd167, 8'd177, 8'd154, 8'd97, 8'd149, 8'd158, 8'd75, 8'd147, 8'd89, 8'd126, 8'd125, 8'd140, 8'd108, 8'd79, 8'd145, 8'd105, 8'd124, 8'd70, 8'd156, 8'd87, 8'd110, 8'd92, 8'd103, 8'd59, 8'd147, 8'd116, 8'd144, 8'd94, 8'd175, 8'd98, 8'd101, 8'd129, 8'd156, 8'd147, 8'd71, 8'd135, 8'd139, 8'd121, 8'd124, 8'd146, 8'd95, 8'd92, 8'd120, 8'd92, 8'd84, 8'd119, 8'd134, 8'd128, 8'd71, 8'd41, 8'd44, 8'd85, 8'd119, 8'd156, 8'd131, 8'd86, 8'd108, 8'd166, 8'd154, 8'd125, 8'd111, 8'd109, 8'd131, 8'd136, 8'd128, 8'd54, 8'd148, 8'd156, 8'd95, 8'd56, 8'd92, 8'd110, 8'd99, 8'd127, 8'd97, 8'd66, 8'd96, 8'd83, 8'd124, 8'd97, 8'd69, 8'd158, 8'd102, 8'd118, 8'd149, 8'd148, 8'd152, 8'd140, 8'd80, 8'd164, 8'd92, 8'd65, 8'd47, 8'd61, 8'd129, 8'd62, 8'd129, 8'd132, 8'd73, 8'd118, 8'd109, 8'd115, 8'd71, 8'd147, 8'd116, 8'd55, 8'd113, 8'd132, 8'd68, 8'd126, 8'd136, 8'd152, 8'd153, 8'd139, 8'd169, 8'd172, 8'd105, 8'd81, 8'd65, 8'd142, 8'd138, 8'd56, 8'd70, 8'd119, 8'd97, 8'd75, 8'd110, 8'd113, 8'd98, 8'd83, 8'd153, 8'd138, 8'd70, 8'd51, 8'd107, 8'd56, 8'd64, 8'd108, 8'd157, 8'd134, 8'd134, 8'd130, 8'd112, 8'd131, 8'd78, 8'd117, 8'd131, 8'd159, 8'd149, 8'd96, 8'd72, 8'd118, 8'd97, 8'd102, 8'd155, 8'd73, 8'd104, 8'd83, 8'd133, 8'd139, 8'd143, 8'd107, 8'd118, 8'd150, 8'd68, 8'd127, 8'd104, 8'd56, 8'd83, 8'd125, 8'd86, 8'd69, 8'd119, 8'd131, 8'd68, 8'd85, 8'd129, 8'd115, 8'd132, 8'd103, 8'd90, 8'd141, 8'd164, 8'd79, 8'd118, 8'd73, 8'd160, 8'd91, 8'd157, 8'd73, 8'd145, 8'd92, 8'd99, 8'd112, 8'd134, 8'd70, 8'd44, 8'd111, 8'd79, 8'd75, 8'd117, 8'd74, 8'd127, 8'd117, 8'd50, 8'd133, 8'd133, 8'd163, 8'd130, 8'd172, 8'd93, 8'd128, 8'd158, 8'd99, 8'd143, 8'd96, 8'd102, 8'd138, 8'd89, 8'd113, 8'd95, 8'd126, 8'd97, 8'd89, 8'd28, 8'd118, 8'd58, 8'd59, 8'd72, 8'd74, 8'd27, 8'd118, 8'd96, 8'd105, 8'd150, 8'd104, 8'd131, 8'd117, 8'd71, 8'd118, 8'd73, 8'd149, 8'd89, 8'd118, 8'd98, 8'd125, 8'd73, 8'd169, 8'd174, 8'd170, 8'd108, 8'd150, 8'd74, 8'd115, 8'd138, 8'd126, 8'd126, 8'd113, 8'd92, 8'd79, 8'd74, 8'd117, 8'd157, 8'd115, 8'd63, 8'd140, 8'd86, 8'd149, 8'd125, 8'd168, 8'd148, 8'd135, 8'd112, 8'd141, 8'd107, 8'd148, 8'd146, 8'd124, 8'd98, 8'd121, 8'd86, 8'd129, 8'd144, 8'd104, 8'd115, 8'd172, 8'd153, 8'd118, 8'd121, 8'd104, 8'd141, 8'd84, 8'd96, 8'd123, 8'd84, 8'd142, 8'd94, 8'd93, 8'd136, 8'd142, 8'd164, 8'd87, 8'd108, 8'd82, 8'd143, 8'd75, 8'd109, 8'd97, 8'd75, 8'd147, 8'd112, 8'd104, 8'd158, 8'd88, 8'd79, 8'd129, 8'd90, 8'd154, 8'd144, 8'd169, 8'd99, 8'd137, 8'd83, 8'd102, 8'd93, 8'd112, 8'd96})
) cell_0_58 (
    .clk(clk),
    .input_index(index_0_57_58),
    .input_value(value_0_57_58),
    .input_result(result_0_57_58),
    .input_enable(enable_0_57_58),
    .output_index(index_0_58_59),
    .output_value(value_0_58_59),
    .output_result(result_0_58_59),
    .output_enable(enable_0_58_59)
);

wire [10-1:0] index_0_59_60;
wire [`DATA_WIDTH-1:0] value_0_59_60;
wire [`DATA_WIDTH*4:0] result_0_59_60;
wire enable_0_59_60;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd120, 8'd152, 8'd141, 8'd167, 8'd145, 8'd108, 8'd79, 8'd145, 8'd122, 8'd137, 8'd39, 8'd57, 8'd96, 8'd140, 8'd138, 8'd105, 8'd73, 8'd120, 8'd149, 8'd157, 8'd78, 8'd124, 8'd159, 8'd98, 8'd99, 8'd139, 8'd122, 8'd144, 8'd154, 8'd168, 8'd123, 8'd104, 8'd161, 8'd91, 8'd88, 8'd144, 8'd136, 8'd113, 8'd139, 8'd124, 8'd104, 8'd175, 8'd189, 8'd99, 8'd141, 8'd155, 8'd148, 8'd123, 8'd171, 8'd183, 8'd114, 8'd126, 8'd108, 8'd156, 8'd132, 8'd97, 8'd158, 8'd66, 8'd83, 8'd127, 8'd167, 8'd140, 8'd178, 8'd175, 8'd137, 8'd176, 8'd129, 8'd156, 8'd115, 8'd124, 8'd133, 8'd129, 8'd112, 8'd141, 8'd108, 8'd153, 8'd97, 8'd168, 8'd106, 8'd89, 8'd66, 8'd142, 8'd112, 8'd132, 8'd144, 8'd128, 8'd93, 8'd157, 8'd126, 8'd128, 8'd118, 8'd145, 8'd105, 8'd149, 8'd139, 8'd150, 8'd153, 8'd75, 8'd85, 8'd120, 8'd158, 8'd168, 8'd146, 8'd86, 8'd142, 8'd165, 8'd123, 8'd143, 8'd115, 8'd112, 8'd130, 8'd170, 8'd155, 8'd140, 8'd108, 8'd168, 8'd111, 8'd132, 8'd90, 8'd104, 8'd115, 8'd87, 8'd152, 8'd92, 8'd63, 8'd148, 8'd124, 8'd120, 8'd145, 8'd152, 8'd149, 8'd154, 8'd124, 8'd77, 8'd112, 8'd68, 8'd88, 8'd57, 8'd109, 8'd131, 8'd119, 8'd157, 8'd140, 8'd118, 8'd105, 8'd169, 8'd114, 8'd125, 8'd138, 8'd121, 8'd90, 8'd84, 8'd157, 8'd144, 8'd76, 8'd87, 8'd148, 8'd112, 8'd113, 8'd116, 8'd77, 8'd59, 8'd75, 8'd94, 8'd143, 8'd70, 8'd150, 8'd148, 8'd126, 8'd66, 8'd126, 8'd102, 8'd178, 8'd113, 8'd160, 8'd127, 8'd92, 8'd85, 8'd132, 8'd160, 8'd156, 8'd93, 8'd99, 8'd74, 8'd81, 8'd108, 8'd116, 8'd113, 8'd77, 8'd95, 8'd99, 8'd137, 8'd61, 8'd139, 8'd120, 8'd73, 8'd106, 8'd73, 8'd158, 8'd93, 8'd102, 8'd139, 8'd141, 8'd144, 8'd84, 8'd83, 8'd127, 8'd129, 8'd63, 8'd94, 8'd144, 8'd55, 8'd63, 8'd139, 8'd145, 8'd79, 8'd152, 8'd68, 8'd127, 8'd86, 8'd61, 8'd119, 8'd143, 8'd102, 8'd113, 8'd131, 8'd82, 8'd79, 8'd86, 8'd102, 8'd151, 8'd83, 8'd116, 8'd144, 8'd134, 8'd88, 8'd98, 8'd137, 8'd70, 8'd134, 8'd102, 8'd58, 8'd104, 8'd103, 8'd76, 8'd171, 8'd81, 8'd65, 8'd70, 8'd78, 8'd85, 8'd155, 8'd87, 8'd131, 8'd113, 8'd164, 8'd98, 8'd89, 8'd132, 8'd150, 8'd117, 8'd136, 8'd81, 8'd167, 8'd177, 8'd86, 8'd129, 8'd129, 8'd124, 8'd81, 8'd117, 8'd143, 8'd165, 8'd125, 8'd131, 8'd80, 8'd57, 8'd101, 8'd137, 8'd143, 8'd87, 8'd67, 8'd109, 8'd131, 8'd110, 8'd124, 8'd144, 8'd106, 8'd107, 8'd147, 8'd144, 8'd91, 8'd83, 8'd83, 8'd106, 8'd130, 8'd122, 8'd162, 8'd75, 8'd125, 8'd118, 8'd97, 8'd104, 8'd64, 8'd95, 8'd89, 8'd72, 8'd89, 8'd158, 8'd102, 8'd110, 8'd73, 8'd143, 8'd141, 8'd78, 8'd127, 8'd93, 8'd151, 8'd100, 8'd181, 8'd127, 8'd58, 8'd121, 8'd118, 8'd84, 8'd112, 8'd113, 8'd92, 8'd134, 8'd155, 8'd151, 8'd125, 8'd147, 8'd51, 8'd104, 8'd143, 8'd150, 8'd130, 8'd133, 8'd75, 8'd54, 8'd152, 8'd138, 8'd167, 8'd100, 8'd131, 8'd179, 8'd120, 8'd139, 8'd135, 8'd85, 8'd78, 8'd91, 8'd160, 8'd143, 8'd107, 8'd150, 8'd116, 8'd87, 8'd171, 8'd115, 8'd63, 8'd77, 8'd137, 8'd79, 8'd93, 8'd42, 8'd104, 8'd118, 8'd101, 8'd170, 8'd152, 8'd83, 8'd118, 8'd163, 8'd126, 8'd160, 8'd152, 8'd147, 8'd126, 8'd136, 8'd182, 8'd84, 8'd108, 8'd139, 8'd126, 8'd185, 8'd123, 8'd92, 8'd58, 8'd107, 8'd85, 8'd74, 8'd73, 8'd75, 8'd13, 8'd96, 8'd95, 8'd114, 8'd120, 8'd158, 8'd158, 8'd126, 8'd165, 8'd148, 8'd134, 8'd152, 8'd173, 8'd130, 8'd93, 8'd147, 8'd139, 8'd120, 8'd109, 8'd186, 8'd152, 8'd147, 8'd105, 8'd143, 8'd145, 8'd125, 8'd132, 8'd66, 8'd31, 8'd63, 8'd110, 8'd154, 8'd128, 8'd125, 8'd143, 8'd156, 8'd97, 8'd71, 8'd61, 8'd84, 8'd128, 8'd141, 8'd173, 8'd84, 8'd105, 8'd133, 8'd105, 8'd122, 8'd137, 8'd144, 8'd108, 8'd100, 8'd143, 8'd145, 8'd125, 8'd87, 8'd146, 8'd117, 8'd77, 8'd114, 8'd159, 8'd147, 8'd143, 8'd155, 8'd123, 8'd99, 8'd137, 8'd150, 8'd163, 8'd155, 8'd113, 8'd152, 8'd167, 8'd126, 8'd179, 8'd132, 8'd62, 8'd97, 8'd91, 8'd133, 8'd152, 8'd145, 8'd173, 8'd119, 8'd176, 8'd79, 8'd102, 8'd161, 8'd76, 8'd136, 8'd119, 8'd110, 8'd133, 8'd88, 8'd63, 8'd135, 8'd78, 8'd124, 8'd130, 8'd114, 8'd155, 8'd111, 8'd157, 8'd151, 8'd73, 8'd134, 8'd111, 8'd144, 8'd98, 8'd150, 8'd179, 8'd188, 8'd134, 8'd105, 8'd108, 8'd126, 8'd154, 8'd127, 8'd83, 8'd81, 8'd144, 8'd154, 8'd80, 8'd113, 8'd89, 8'd108, 8'd175, 8'd82, 8'd157, 8'd129, 8'd156, 8'd86, 8'd117, 8'd99, 8'd102, 8'd55, 8'd92, 8'd136, 8'd93, 8'd104, 8'd137, 8'd162, 8'd100, 8'd74, 8'd72, 8'd86, 8'd89, 8'd103, 8'd141, 8'd164, 8'd126, 8'd99, 8'd91, 8'd92, 8'd119, 8'd135, 8'd102, 8'd146, 8'd105, 8'd43, 8'd52, 8'd110, 8'd142, 8'd82, 8'd129, 8'd136, 8'd162, 8'd155, 8'd102, 8'd61, 8'd88, 8'd81, 8'd146, 8'd95, 8'd134, 8'd178, 8'd152, 8'd115, 8'd139, 8'd171, 8'd156, 8'd107, 8'd104, 8'd79, 8'd104, 8'd129, 8'd109, 8'd36, 8'd107, 8'd65, 8'd143, 8'd117, 8'd117, 8'd154, 8'd181, 8'd150, 8'd169, 8'd124, 8'd78, 8'd88, 8'd131, 8'd77, 8'd83, 8'd111, 8'd179, 8'd170, 8'd179, 8'd151, 8'd91, 8'd120, 8'd113, 8'd113, 8'd149, 8'd56, 8'd75, 8'd60, 8'd108, 8'd146, 8'd89, 8'd78, 8'd75, 8'd157, 8'd111, 8'd89, 8'd171, 8'd74, 8'd75, 8'd148, 8'd83, 8'd103, 8'd94, 8'd146, 8'd91, 8'd136, 8'd116, 8'd118, 8'd173, 8'd131, 8'd77, 8'd64, 8'd83, 8'd150, 8'd51, 8'd135, 8'd51, 8'd146, 8'd144, 8'd101, 8'd136, 8'd125, 8'd86, 8'd137, 8'd103, 8'd147, 8'd85, 8'd94, 8'd64, 8'd107, 8'd77, 8'd90, 8'd135, 8'd96, 8'd50, 8'd136, 8'd88, 8'd95, 8'd118, 8'd62, 8'd138, 8'd134, 8'd80, 8'd75, 8'd139, 8'd70, 8'd107, 8'd74, 8'd71, 8'd150, 8'd91, 8'd133, 8'd159, 8'd67, 8'd154, 8'd139, 8'd105, 8'd149, 8'd102, 8'd119, 8'd60, 8'd56, 8'd74, 8'd39, 8'd88, 8'd137, 8'd140, 8'd138, 8'd59, 8'd122, 8'd86, 8'd121, 8'd129, 8'd90, 8'd107, 8'd91, 8'd72, 8'd152, 8'd137, 8'd80, 8'd148, 8'd55, 8'd70, 8'd89, 8'd139, 8'd60, 8'd53, 8'd93, 8'd66, 8'd42, 8'd120, 8'd67, 8'd62, 8'd119, 8'd99, 8'd47, 8'd88, 8'd84, 8'd136, 8'd97, 8'd96, 8'd140, 8'd75, 8'd155, 8'd117, 8'd79, 8'd95, 8'd98, 8'd113, 8'd152, 8'd136, 8'd128, 8'd115, 8'd117, 8'd79, 8'd100, 8'd130, 8'd116, 8'd124, 8'd99, 8'd83, 8'd62, 8'd123, 8'd123, 8'd67, 8'd70, 8'd124, 8'd81, 8'd117, 8'd138, 8'd97, 8'd113, 8'd166, 8'd105, 8'd115, 8'd74, 8'd147, 8'd155, 8'd125, 8'd81, 8'd122, 8'd95, 8'd78, 8'd167, 8'd154, 8'd139, 8'd130, 8'd72, 8'd139, 8'd77, 8'd70, 8'd143, 8'd83, 8'd80, 8'd86, 8'd108, 8'd79, 8'd97, 8'd166, 8'd120, 8'd144})
) cell_0_59 (
    .clk(clk),
    .input_index(index_0_58_59),
    .input_value(value_0_58_59),
    .input_result(result_0_58_59),
    .input_enable(enable_0_58_59),
    .output_index(index_0_59_60),
    .output_value(value_0_59_60),
    .output_result(result_0_59_60),
    .output_enable(enable_0_59_60)
);

wire [10-1:0] index_0_60_61;
wire [`DATA_WIDTH-1:0] value_0_60_61;
wire [`DATA_WIDTH*4:0] result_0_60_61;
wire enable_0_60_61;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd133, 8'd144, 8'd131, 8'd85, 8'd60, 8'd148, 8'd86, 8'd105, 8'd73, 8'd73, 8'd69, 8'd70, 8'd147, 8'd79, 8'd134, 8'd82, 8'd70, 8'd83, 8'd65, 8'd131, 8'd79, 8'd69, 8'd114, 8'd75, 8'd82, 8'd165, 8'd155, 8'd148, 8'd164, 8'd93, 8'd110, 8'd119, 8'd112, 8'd86, 8'd105, 8'd127, 8'd84, 8'd114, 8'd140, 8'd95, 8'd86, 8'd79, 8'd132, 8'd94, 8'd108, 8'd161, 8'd79, 8'd152, 8'd86, 8'd141, 8'd100, 8'd91, 8'd105, 8'd122, 8'd145, 8'd88, 8'd101, 8'd112, 8'd98, 8'd88, 8'd130, 8'd101, 8'd137, 8'd188, 8'd117, 8'd145, 8'd130, 8'd76, 8'd88, 8'd61, 8'd146, 8'd71, 8'd117, 8'd62, 8'd124, 8'd76, 8'd157, 8'd127, 8'd169, 8'd70, 8'd126, 8'd136, 8'd126, 8'd157, 8'd80, 8'd78, 8'd85, 8'd68, 8'd129, 8'd169, 8'd114, 8'd92, 8'd170, 8'd137, 8'd156, 8'd92, 8'd121, 8'd73, 8'd104, 8'd134, 8'd122, 8'd132, 8'd141, 8'd73, 8'd126, 8'd72, 8'd119, 8'd96, 8'd106, 8'd139, 8'd79, 8'd95, 8'd114, 8'd138, 8'd135, 8'd157, 8'd108, 8'd156, 8'd160, 8'd115, 8'd82, 8'd74, 8'd105, 8'd143, 8'd93, 8'd75, 8'd48, 8'd112, 8'd88, 8'd143, 8'd155, 8'd99, 8'd104, 8'd131, 8'd133, 8'd57, 8'd149, 8'd91, 8'd90, 8'd101, 8'd171, 8'd156, 8'd72, 8'd86, 8'd166, 8'd158, 8'd116, 8'd147, 8'd127, 8'd139, 8'd169, 8'd83, 8'd78, 8'd66, 8'd141, 8'd109, 8'd145, 8'd74, 8'd64, 8'd156, 8'd71, 8'd86, 8'd154, 8'd145, 8'd125, 8'd137, 8'd168, 8'd122, 8'd172, 8'd84, 8'd79, 8'd115, 8'd105, 8'd65, 8'd143, 8'd86, 8'd144, 8'd121, 8'd86, 8'd148, 8'd103, 8'd64, 8'd64, 8'd62, 8'd90, 8'd120, 8'd131, 8'd94, 8'd89, 8'd74, 8'd173, 8'd73, 8'd100, 8'd90, 8'd154, 8'd113, 8'd162, 8'd73, 8'd115, 8'd58, 8'd98, 8'd136, 8'd120, 8'd106, 8'd77, 8'd161, 8'd69, 8'd164, 8'd76, 8'd60, 8'd83, 8'd95, 8'd113, 8'd92, 8'd125, 8'd148, 8'd67, 8'd108, 8'd161, 8'd135, 8'd152, 8'd124, 8'd140, 8'd143, 8'd114, 8'd134, 8'd87, 8'd77, 8'd98, 8'd105, 8'd107, 8'd93, 8'd114, 8'd103, 8'd111, 8'd162, 8'd141, 8'd84, 8'd95, 8'd116, 8'd121, 8'd91, 8'd68, 8'd151, 8'd133, 8'd151, 8'd138, 8'd65, 8'd78, 8'd119, 8'd155, 8'd155, 8'd130, 8'd71, 8'd87, 8'd34, 8'd58, 8'd130, 8'd87, 8'd125, 8'd142, 8'd146, 8'd67, 8'd149, 8'd68, 8'd153, 8'd130, 8'd102, 8'd91, 8'd139, 8'd78, 8'd141, 8'd131, 8'd127, 8'd85, 8'd105, 8'd119, 8'd111, 8'd125, 8'd142, 8'd70, 8'd68, 8'd46, 8'd36, 8'd87, 8'd138, 8'd81, 8'd60, 8'd82, 8'd74, 8'd107, 8'd116, 8'd119, 8'd72, 8'd116, 8'd95, 8'd145, 8'd145, 8'd130, 8'd110, 8'd167, 8'd62, 8'd70, 8'd114, 8'd96, 8'd102, 8'd94, 8'd121, 8'd98, 8'd45, 8'd43, 8'd108, 8'd125, 8'd129, 8'd92, 8'd137, 8'd92, 8'd142, 8'd51, 8'd98, 8'd121, 8'd66, 8'd147, 8'd139, 8'd146, 8'd147, 8'd102, 8'd146, 8'd136, 8'd122, 8'd94, 8'd127, 8'd102, 8'd126, 8'd81, 8'd133, 8'd138, 8'd108, 8'd111, 8'd105, 8'd101, 8'd119, 8'd134, 8'd78, 8'd145, 8'd56, 8'd133, 8'd118, 8'd83, 8'd104, 8'd139, 8'd129, 8'd140, 8'd116, 8'd110, 8'd165, 8'd110, 8'd120, 8'd99, 8'd139, 8'd141, 8'd112, 8'd79, 8'd131, 8'd138, 8'd54, 8'd97, 8'd124, 8'd88, 8'd166, 8'd100, 8'd134, 8'd64, 8'd123, 8'd84, 8'd112, 8'd127, 8'd92, 8'd188, 8'd178, 8'd135, 8'd107, 8'd104, 8'd184, 8'd128, 8'd172, 8'd118, 8'd85, 8'd74, 8'd73, 8'd101, 8'd121, 8'd132, 8'd80, 8'd58, 8'd95, 8'd133, 8'd89, 8'd162, 8'd81, 8'd122, 8'd154, 8'd158, 8'd88, 8'd107, 8'd193, 8'd206, 8'd134, 8'd175, 8'd118, 8'd125, 8'd159, 8'd124, 8'd192, 8'd190, 8'd99, 8'd129, 8'd136, 8'd111, 8'd138, 8'd124, 8'd51, 8'd55, 8'd68, 8'd148, 8'd166, 8'd98, 8'd116, 8'd120, 8'd96, 8'd88, 8'd80, 8'd160, 8'd212, 8'd158, 8'd121, 8'd124, 8'd111, 8'd146, 8'd89, 8'd136, 8'd132, 8'd102, 8'd73, 8'd78, 8'd68, 8'd67, 8'd155, 8'd123, 8'd50, 8'd39, 8'd83, 8'd133, 8'd136, 8'd105, 8'd108, 8'd120, 8'd125, 8'd126, 8'd124, 8'd130, 8'd138, 8'd128, 8'd92, 8'd140, 8'd90, 8'd145, 8'd114, 8'd138, 8'd118, 8'd126, 8'd115, 8'd44, 8'd61, 8'd93, 8'd142, 8'd115, 8'd103, 8'd89, 8'd122, 8'd86, 8'd119, 8'd51, 8'd50, 8'd112, 8'd135, 8'd53, 8'd144, 8'd160, 8'd131, 8'd160, 8'd176, 8'd120, 8'd154, 8'd98, 8'd120, 8'd148, 8'd124, 8'd76, 8'd130, 8'd52, 8'd63, 8'd78, 8'd70, 8'd146, 8'd86, 8'd101, 8'd88, 8'd116, 8'd103, 8'd116, 8'd116, 8'd124, 8'd86, 8'd59, 8'd144, 8'd71, 8'd96, 8'd130, 8'd62, 8'd86, 8'd61, 8'd79, 8'd55, 8'd84, 8'd54, 8'd79, 8'd68, 8'd92, 8'd55, 8'd141, 8'd66, 8'd154, 8'd99, 8'd119, 8'd114, 8'd58, 8'd51, 8'd141, 8'd132, 8'd78, 8'd107, 8'd77, 8'd120, 8'd72, 8'd70, 8'd132, 8'd101, 8'd65, 8'd31, 8'd87, 8'd89, 8'd94, 8'd119, 8'd115, 8'd94, 8'd52, 8'd73, 8'd142, 8'd109, 8'd67, 8'd72, 8'd46, 8'd92, 8'd79, 8'd127, 8'd151, 8'd135, 8'd73, 8'd95, 8'd81, 8'd107, 8'd94, 8'd116, 8'd113, 8'd107, 8'd43, 8'd55, 8'd67, 8'd28, 8'd68, 8'd79, 8'd33, 8'd115, 8'd52, 8'd106, 8'd64, 8'd112, 8'd112, 8'd132, 8'd67, 8'd95, 8'd165, 8'd121, 8'd152, 8'd154, 8'd120, 8'd148, 8'd130, 8'd97, 8'd146, 8'd146, 8'd134, 8'd113, 8'd48, 8'd39, 8'd39, 8'd90, 8'd103, 8'd86, 8'd93, 8'd78, 8'd101, 8'd103, 8'd141, 8'd130, 8'd124, 8'd88, 8'd117, 8'd156, 8'd204, 8'd194, 8'd183, 8'd116, 8'd149, 8'd113, 8'd137, 8'd60, 8'd133, 8'd93, 8'd96, 8'd100, 8'd152, 8'd77, 8'd95, 8'd71, 8'd98, 8'd92, 8'd131, 8'd113, 8'd99, 8'd76, 8'd130, 8'd92, 8'd93, 8'd155, 8'd118, 8'd113, 8'd188, 8'd202, 8'd114, 8'd101, 8'd162, 8'd157, 8'd73, 8'd100, 8'd128, 8'd96, 8'd71, 8'd139, 8'd111, 8'd50, 8'd121, 8'd140, 8'd117, 8'd90, 8'd94, 8'd120, 8'd72, 8'd127, 8'd143, 8'd122, 8'd147, 8'd138, 8'd95, 8'd157, 8'd179, 8'd99, 8'd96, 8'd146, 8'd124, 8'd132, 8'd46, 8'd43, 8'd123, 8'd133, 8'd68, 8'd37, 8'd38, 8'd111, 8'd66, 8'd114, 8'd84, 8'd142, 8'd119, 8'd136, 8'd156, 8'd122, 8'd94, 8'd161, 8'd160, 8'd118, 8'd145, 8'd79, 8'd123, 8'd114, 8'd123, 8'd83, 8'd60, 8'd98, 8'd100, 8'd92, 8'd114, 8'd64, 8'd142, 8'd53, 8'd53, 8'd98, 8'd59, 8'd123, 8'd97, 8'd68, 8'd123, 8'd147, 8'd162, 8'd108, 8'd141, 8'd115, 8'd73, 8'd74, 8'd80, 8'd99, 8'd94, 8'd63, 8'd85, 8'd111, 8'd110, 8'd119, 8'd76, 8'd94, 8'd90, 8'd157, 8'd89, 8'd154, 8'd94, 8'd114, 8'd167, 8'd84, 8'd102, 8'd93, 8'd147, 8'd135, 8'd112, 8'd78, 8'd147, 8'd125, 8'd151, 8'd128, 8'd75, 8'd123, 8'd151, 8'd90, 8'd86, 8'd159, 8'd120, 8'd133, 8'd139, 8'd87, 8'd159, 8'd133, 8'd72, 8'd131, 8'd148, 8'd99, 8'd104, 8'd104, 8'd73, 8'd147, 8'd84, 8'd122, 8'd128, 8'd117, 8'd153, 8'd94})
) cell_0_60 (
    .clk(clk),
    .input_index(index_0_59_60),
    .input_value(value_0_59_60),
    .input_result(result_0_59_60),
    .input_enable(enable_0_59_60),
    .output_index(index_0_60_61),
    .output_value(value_0_60_61),
    .output_result(result_0_60_61),
    .output_enable(enable_0_60_61)
);

wire [10-1:0] index_0_61_62;
wire [`DATA_WIDTH-1:0] value_0_61_62;
wire [`DATA_WIDTH*4:0] result_0_61_62;
wire enable_0_61_62;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd160, 8'd84, 8'd120, 8'd126, 8'd85, 8'd145, 8'd69, 8'd134, 8'd64, 8'd79, 8'd137, 8'd110, 8'd119, 8'd118, 8'd63, 8'd128, 8'd131, 8'd130, 8'd95, 8'd73, 8'd70, 8'd102, 8'd140, 8'd86, 8'd95, 8'd168, 8'd129, 8'd83, 8'd94, 8'd86, 8'd73, 8'd81, 8'd116, 8'd83, 8'd113, 8'd148, 8'd100, 8'd86, 8'd116, 8'd83, 8'd121, 8'd196, 8'd152, 8'd181, 8'd99, 8'd121, 8'd165, 8'd97, 8'd178, 8'd103, 8'd191, 8'd136, 8'd102, 8'd105, 8'd156, 8'd93, 8'd156, 8'd156, 8'd81, 8'd109, 8'd170, 8'd180, 8'd109, 8'd115, 8'd180, 8'd133, 8'd161, 8'd154, 8'd138, 8'd108, 8'd93, 8'd108, 8'd158, 8'd100, 8'd100, 8'd97, 8'd181, 8'd177, 8'd168, 8'd100, 8'd160, 8'd139, 8'd166, 8'd132, 8'd129, 8'd73, 8'd157, 8'd133, 8'd126, 8'd96, 8'd175, 8'd149, 8'd165, 8'd97, 8'd84, 8'd158, 8'd145, 8'd90, 8'd98, 8'd70, 8'd91, 8'd165, 8'd153, 8'd135, 8'd186, 8'd162, 8'd166, 8'd125, 8'd136, 8'd151, 8'd73, 8'd109, 8'd140, 8'd101, 8'd135, 8'd110, 8'd119, 8'd157, 8'd149, 8'd104, 8'd105, 8'd82, 8'd74, 8'd112, 8'd71, 8'd53, 8'd113, 8'd88, 8'd125, 8'd86, 8'd151, 8'd156, 8'd107, 8'd156, 8'd151, 8'd130, 8'd105, 8'd124, 8'd127, 8'd130, 8'd91, 8'd156, 8'd138, 8'd140, 8'd85, 8'd114, 8'd139, 8'd165, 8'd130, 8'd70, 8'd133, 8'd72, 8'd144, 8'd153, 8'd61, 8'd125, 8'd92, 8'd64, 8'd124, 8'd124, 8'd116, 8'd58, 8'd121, 8'd85, 8'd93, 8'd84, 8'd96, 8'd157, 8'd158, 8'd82, 8'd126, 8'd147, 8'd140, 8'd81, 8'd161, 8'd95, 8'd109, 8'd113, 8'd131, 8'd126, 8'd125, 8'd113, 8'd152, 8'd130, 8'd73, 8'd91, 8'd103, 8'd64, 8'd115, 8'd68, 8'd91, 8'd70, 8'd71, 8'd76, 8'd137, 8'd119, 8'd84, 8'd102, 8'd158, 8'd97, 8'd134, 8'd102, 8'd78, 8'd147, 8'd141, 8'd100, 8'd114, 8'd142, 8'd73, 8'd118, 8'd100, 8'd117, 8'd77, 8'd92, 8'd136, 8'd115, 8'd81, 8'd98, 8'd100, 8'd140, 8'd115, 8'd158, 8'd113, 8'd150, 8'd157, 8'd183, 8'd78, 8'd73, 8'd103, 8'd59, 8'd58, 8'd125, 8'd152, 8'd134, 8'd84, 8'd108, 8'd156, 8'd137, 8'd76, 8'd62, 8'd132, 8'd125, 8'd72, 8'd110, 8'd56, 8'd87, 8'd123, 8'd46, 8'd104, 8'd132, 8'd88, 8'd107, 8'd116, 8'd176, 8'd101, 8'd63, 8'd109, 8'd83, 8'd129, 8'd163, 8'd82, 8'd114, 8'd70, 8'd76, 8'd176, 8'd125, 8'd94, 8'd101, 8'd133, 8'd80, 8'd141, 8'd98, 8'd62, 8'd148, 8'd134, 8'd132, 8'd81, 8'd100, 8'd132, 8'd136, 8'd104, 8'd162, 8'd129, 8'd131, 8'd143, 8'd140, 8'd86, 8'd101, 8'd83, 8'd94, 8'd142, 8'd154, 8'd172, 8'd101, 8'd158, 8'd151, 8'd134, 8'd87, 8'd109, 8'd75, 8'd160, 8'd119, 8'd80, 8'd126, 8'd121, 8'd146, 8'd154, 8'd144, 8'd154, 8'd133, 8'd96, 8'd96, 8'd100, 8'd127, 8'd119, 8'd139, 8'd137, 8'd148, 8'd104, 8'd139, 8'd116, 8'd166, 8'd83, 8'd78, 8'd139, 8'd103, 8'd143, 8'd141, 8'd83, 8'd119, 8'd137, 8'd77, 8'd126, 8'd118, 8'd140, 8'd150, 8'd155, 8'd171, 8'd59, 8'd61, 8'd94, 8'd103, 8'd148, 8'd79, 8'd172, 8'd122, 8'd135, 8'd183, 8'd135, 8'd87, 8'd154, 8'd96, 8'd136, 8'd103, 8'd166, 8'd161, 8'd85, 8'd97, 8'd152, 8'd138, 8'd151, 8'd85, 8'd148, 8'd156, 8'd148, 8'd62, 8'd103, 8'd122, 8'd63, 8'd110, 8'd92, 8'd94, 8'd163, 8'd166, 8'd179, 8'd127, 8'd159, 8'd140, 8'd151, 8'd150, 8'd83, 8'd168, 8'd144, 8'd145, 8'd132, 8'd96, 8'd115, 8'd174, 8'd145, 8'd135, 8'd117, 8'd112, 8'd89, 8'd78, 8'd140, 8'd45, 8'd134, 8'd139, 8'd154, 8'd166, 8'd165, 8'd127, 8'd112, 8'd145, 8'd183, 8'd159, 8'd110, 8'd126, 8'd135, 8'd117, 8'd180, 8'd149, 8'd172, 8'd151, 8'd163, 8'd160, 8'd80, 8'd96, 8'd140, 8'd152, 8'd62, 8'd135, 8'd71, 8'd132, 8'd98, 8'd136, 8'd172, 8'd146, 8'd117, 8'd100, 8'd107, 8'd121, 8'd126, 8'd118, 8'd90, 8'd91, 8'd114, 8'd140, 8'd119, 8'd133, 8'd162, 8'd166, 8'd83, 8'd151, 8'd77, 8'd139, 8'd85, 8'd87, 8'd112, 8'd135, 8'd97, 8'd100, 8'd56, 8'd65, 8'd91, 8'd97, 8'd104, 8'd93, 8'd98, 8'd123, 8'd99, 8'd133, 8'd52, 8'd154, 8'd80, 8'd131, 8'd155, 8'd165, 8'd114, 8'd126, 8'd86, 8'd118, 8'd126, 8'd108, 8'd81, 8'd103, 8'd61, 8'd55, 8'd109, 8'd58, 8'd82, 8'd69, 8'd67, 8'd58, 8'd110, 8'd153, 8'd116, 8'd155, 8'd144, 8'd135, 8'd77, 8'd163, 8'd101, 8'd127, 8'd129, 8'd122, 8'd91, 8'd130, 8'd142, 8'd111, 8'd48, 8'd68, 8'd88, 8'd131, 8'd88, 8'd76, 8'd83, 8'd46, 8'd64, 8'd76, 8'd71, 8'd59, 8'd142, 8'd62, 8'd81, 8'd68, 8'd135, 8'd108, 8'd95, 8'd129, 8'd160, 8'd115, 8'd78, 8'd93, 8'd99, 8'd115, 8'd74, 8'd68, 8'd114, 8'd97, 8'd86, 8'd124, 8'd81, 8'd63, 8'd65, 8'd42, 8'd31, 8'd92, 8'd129, 8'd151, 8'd127, 8'd69, 8'd152, 8'd156, 8'd158, 8'd121, 8'd99, 8'd121, 8'd125, 8'd123, 8'd150, 8'd160, 8'd117, 8'd60, 8'd113, 8'd74, 8'd63, 8'd85, 8'd86, 8'd115, 8'd79, 8'd109, 8'd58, 8'd98, 8'd88, 8'd96, 8'd113, 8'd123, 8'd128, 8'd117, 8'd124, 8'd172, 8'd126, 8'd141, 8'd131, 8'd128, 8'd134, 8'd113, 8'd135, 8'd142, 8'd82, 8'd108, 8'd132, 8'd142, 8'd138, 8'd121, 8'd74, 8'd75, 8'd113, 8'd153, 8'd81, 8'd62, 8'd60, 8'd114, 8'd117, 8'd149, 8'd108, 8'd107, 8'd92, 8'd137, 8'd130, 8'd149, 8'd101, 8'd85, 8'd84, 8'd121, 8'd129, 8'd103, 8'd136, 8'd81, 8'd149, 8'd167, 8'd132, 8'd97, 8'd150, 8'd96, 8'd165, 8'd93, 8'd125, 8'd102, 8'd144, 8'd144, 8'd140, 8'd60, 8'd87, 8'd83, 8'd91, 8'd100, 8'd123, 8'd144, 8'd145, 8'd74, 8'd114, 8'd122, 8'd90, 8'd155, 8'd115, 8'd92, 8'd103, 8'd168, 8'd94, 8'd97, 8'd120, 8'd77, 8'd157, 8'd118, 8'd116, 8'd88, 8'd168, 8'd138, 8'd116, 8'd182, 8'd125, 8'd104, 8'd115, 8'd75, 8'd48, 8'd80, 8'd96, 8'd85, 8'd82, 8'd67, 8'd126, 8'd99, 8'd99, 8'd90, 8'd92, 8'd114, 8'd65, 8'd87, 8'd107, 8'd108, 8'd120, 8'd116, 8'd109, 8'd128, 8'd96, 8'd156, 8'd127, 8'd146, 8'd88, 8'd152, 8'd72, 8'd90, 8'd64, 8'd45, 8'd68, 8'd82, 8'd69, 8'd104, 8'd147, 8'd93, 8'd138, 8'd147, 8'd100, 8'd72, 8'd155, 8'd97, 8'd136, 8'd129, 8'd167, 8'd121, 8'd123, 8'd112, 8'd122, 8'd90, 8'd136, 8'd110, 8'd104, 8'd81, 8'd133, 8'd124, 8'd90, 8'd71, 8'd57, 8'd109, 8'd95, 8'd106, 8'd69, 8'd137, 8'd122, 8'd108, 8'd68, 8'd128, 8'd101, 8'd108, 8'd121, 8'd159, 8'd109, 8'd130, 8'd109, 8'd158, 8'd61, 8'd74, 8'd72, 8'd102, 8'd135, 8'd150, 8'd146, 8'd81, 8'd135, 8'd149, 8'd94, 8'd51, 8'd132, 8'd70, 8'd126, 8'd149, 8'd64, 8'd145, 8'd95, 8'd158, 8'd104, 8'd161, 8'd102, 8'd130, 8'd90, 8'd76, 8'd130, 8'd136, 8'd92, 8'd106, 8'd145, 8'd160, 8'd95, 8'd159, 8'd103, 8'd156, 8'd81, 8'd154, 8'd64, 8'd119, 8'd150, 8'd148, 8'd162, 8'd115, 8'd116, 8'd144, 8'd112, 8'd92, 8'd118, 8'd93, 8'd82, 8'd144})
) cell_0_61 (
    .clk(clk),
    .input_index(index_0_60_61),
    .input_value(value_0_60_61),
    .input_result(result_0_60_61),
    .input_enable(enable_0_60_61),
    .output_index(index_0_61_62),
    .output_value(value_0_61_62),
    .output_result(result_0_61_62),
    .output_enable(enable_0_61_62)
);

wire [10-1:0] index_0_62_63;
wire [`DATA_WIDTH-1:0] value_0_62_63;
wire [`DATA_WIDTH*4:0] result_0_62_63;
wire enable_0_62_63;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd100, 8'd87, 8'd142, 8'd113, 8'd62, 8'd122, 8'd113, 8'd108, 8'd106, 8'd162, 8'd88, 8'd130, 8'd152, 8'd128, 8'd61, 8'd108, 8'd126, 8'd144, 8'd129, 8'd154, 8'd155, 8'd102, 8'd127, 8'd144, 8'd94, 8'd158, 8'd79, 8'd161, 8'd82, 8'd162, 8'd151, 8'd105, 8'd149, 8'd166, 8'd165, 8'd180, 8'd107, 8'd147, 8'd128, 8'd125, 8'd177, 8'd121, 8'd188, 8'd134, 8'd180, 8'd167, 8'd122, 8'd181, 8'd105, 8'd182, 8'd112, 8'd113, 8'd143, 8'd163, 8'd103, 8'd88, 8'd169, 8'd108, 8'd78, 8'd138, 8'd162, 8'd91, 8'd111, 8'd143, 8'd169, 8'd111, 8'd161, 8'd117, 8'd123, 8'd88, 8'd153, 8'd80, 8'd105, 8'd110, 8'd143, 8'd123, 8'd174, 8'd165, 8'd132, 8'd169, 8'd162, 8'd155, 8'd169, 8'd111, 8'd142, 8'd75, 8'd157, 8'd111, 8'd117, 8'd167, 8'd158, 8'd129, 8'd137, 8'd71, 8'd78, 8'd87, 8'd91, 8'd147, 8'd98, 8'd142, 8'd130, 8'd97, 8'd83, 8'd113, 8'd97, 8'd75, 8'd162, 8'd118, 8'd151, 8'd143, 8'd143, 8'd110, 8'd88, 8'd109, 8'd171, 8'd109, 8'd158, 8'd159, 8'd186, 8'd104, 8'd146, 8'd78, 8'd76, 8'd106, 8'd67, 8'd94, 8'd96, 8'd120, 8'd81, 8'd123, 8'd148, 8'd132, 8'd136, 8'd111, 8'd95, 8'd63, 8'd74, 8'd142, 8'd157, 8'd158, 8'd152, 8'd152, 8'd171, 8'd162, 8'd111, 8'd187, 8'd175, 8'd137, 8'd141, 8'd78, 8'd103, 8'd88, 8'd92, 8'd121, 8'd102, 8'd124, 8'd174, 8'd81, 8'd104, 8'd102, 8'd151, 8'd127, 8'd114, 8'd104, 8'd69, 8'd78, 8'd85, 8'd129, 8'd85, 8'd114, 8'd91, 8'd185, 8'd162, 8'd115, 8'd121, 8'd150, 8'd94, 8'd148, 8'd114, 8'd76, 8'd84, 8'd139, 8'd136, 8'd159, 8'd152, 8'd129, 8'd71, 8'd133, 8'd135, 8'd126, 8'd102, 8'd129, 8'd72, 8'd161, 8'd129, 8'd122, 8'd69, 8'd166, 8'd176, 8'd193, 8'd96, 8'd167, 8'd96, 8'd64, 8'd99, 8'd77, 8'd62, 8'd154, 8'd154, 8'd135, 8'd97, 8'd159, 8'd127, 8'd145, 8'd89, 8'd124, 8'd104, 8'd90, 8'd111, 8'd70, 8'd61, 8'd168, 8'd94, 8'd145, 8'd121, 8'd86, 8'd179, 8'd118, 8'd150, 8'd98, 8'd72, 8'd102, 8'd148, 8'd113, 8'd79, 8'd125, 8'd143, 8'd108, 8'd123, 8'd148, 8'd126, 8'd105, 8'd150, 8'd122, 8'd166, 8'd164, 8'd112, 8'd100, 8'd122, 8'd67, 8'd81, 8'd83, 8'd88, 8'd155, 8'd176, 8'd156, 8'd83, 8'd69, 8'd107, 8'd158, 8'd138, 8'd126, 8'd119, 8'd112, 8'd133, 8'd109, 8'd126, 8'd112, 8'd111, 8'd159, 8'd89, 8'd160, 8'd172, 8'd171, 8'd169, 8'd151, 8'd119, 8'd100, 8'd96, 8'd166, 8'd142, 8'd173, 8'd155, 8'd181, 8'd142, 8'd82, 8'd77, 8'd99, 8'd97, 8'd171, 8'd150, 8'd126, 8'd162, 8'd128, 8'd81, 8'd122, 8'd95, 8'd123, 8'd172, 8'd129, 8'd131, 8'd174, 8'd129, 8'd67, 8'd85, 8'd70, 8'd73, 8'd134, 8'd92, 8'd168, 8'd160, 8'd97, 8'd69, 8'd112, 8'd74, 8'd113, 8'd133, 8'd146, 8'd188, 8'd114, 8'd132, 8'd48, 8'd79, 8'd103, 8'd125, 8'd109, 8'd116, 8'd129, 8'd89, 8'd185, 8'd162, 8'd152, 8'd103, 8'd148, 8'd105, 8'd99, 8'd152, 8'd175, 8'd121, 8'd154, 8'd100, 8'd139, 8'd131, 8'd126, 8'd124, 8'd148, 8'd173, 8'd168, 8'd127, 8'd82, 8'd102, 8'd135, 8'd155, 8'd125, 8'd177, 8'd166, 8'd151, 8'd183, 8'd104, 8'd127, 8'd62, 8'd95, 8'd76, 8'd122, 8'd121, 8'd198, 8'd171, 8'd133, 8'd83, 8'd133, 8'd130, 8'd132, 8'd151, 8'd176, 8'd168, 8'd118, 8'd67, 8'd51, 8'd125, 8'd85, 8'd140, 8'd141, 8'd112, 8'd132, 8'd114, 8'd130, 8'd162, 8'd85, 8'd106, 8'd93, 8'd140, 8'd149, 8'd121, 8'd130, 8'd100, 8'd58, 8'd73, 8'd147, 8'd125, 8'd117, 8'd150, 8'd85, 8'd117, 8'd97, 8'd64, 8'd119, 8'd66, 8'd100, 8'd103, 8'd104, 8'd130, 8'd87, 8'd108, 8'd138, 8'd150, 8'd132, 8'd161, 8'd55, 8'd147, 8'd82, 8'd134, 8'd119, 8'd116, 8'd112, 8'd79, 8'd74, 8'd108, 8'd97, 8'd135, 8'd83, 8'd109, 8'd73, 8'd134, 8'd111, 8'd143, 8'd59, 8'd155, 8'd153, 8'd82, 8'd164, 8'd74, 8'd159, 8'd82, 8'd110, 8'd151, 8'd118, 8'd125, 8'd109, 8'd103, 8'd77, 8'd112, 8'd147, 8'd96, 8'd142, 8'd106, 8'd129, 8'd125, 8'd129, 8'd132, 8'd157, 8'd56, 8'd74, 8'd78, 8'd155, 8'd165, 8'd94, 8'd177, 8'd153, 8'd107, 8'd176, 8'd123, 8'd132, 8'd131, 8'd51, 8'd80, 8'd131, 8'd143, 8'd138, 8'd169, 8'd192, 8'd128, 8'd156, 8'd151, 8'd175, 8'd152, 8'd154, 8'd139, 8'd152, 8'd141, 8'd64, 8'd71, 8'd96, 8'd128, 8'd112, 8'd183, 8'd93, 8'd124, 8'd148, 8'd118, 8'd147, 8'd59, 8'd124, 8'd96, 8'd123, 8'd174, 8'd147, 8'd105, 8'd121, 8'd104, 8'd83, 8'd103, 8'd125, 8'd144, 8'd159, 8'd134, 8'd134, 8'd165, 8'd103, 8'd105, 8'd178, 8'd174, 8'd107, 8'd168, 8'd166, 8'd80, 8'd120, 8'd149, 8'd80, 8'd111, 8'd141, 8'd118, 8'd153, 8'd72, 8'd158, 8'd109, 8'd139, 8'd110, 8'd136, 8'd88, 8'd141, 8'd111, 8'd95, 8'd121, 8'd127, 8'd157, 8'd90, 8'd141, 8'd153, 8'd133, 8'd101, 8'd132, 8'd164, 8'd123, 8'd159, 8'd121, 8'd78, 8'd87, 8'd101, 8'd120, 8'd135, 8'd77, 8'd105, 8'd172, 8'd172, 8'd119, 8'd94, 8'd124, 8'd146, 8'd80, 8'd106, 8'd94, 8'd121, 8'd118, 8'd140, 8'd171, 8'd127, 8'd164, 8'd172, 8'd111, 8'd138, 8'd128, 8'd137, 8'd84, 8'd114, 8'd110, 8'd97, 8'd159, 8'd81, 8'd105, 8'd153, 8'd112, 8'd101, 8'd138, 8'd109, 8'd140, 8'd132, 8'd168, 8'd147, 8'd146, 8'd133, 8'd107, 8'd128, 8'd156, 8'd102, 8'd164, 8'd168, 8'd162, 8'd138, 8'd137, 8'd99, 8'd85, 8'd75, 8'd65, 8'd109, 8'd110, 8'd83, 8'd163, 8'd165, 8'd124, 8'd70, 8'd127, 8'd102, 8'd119, 8'd76, 8'd99, 8'd104, 8'd113, 8'd97, 8'd88, 8'd128, 8'd103, 8'd130, 8'd151, 8'd104, 8'd129, 8'd77, 8'd154, 8'd104, 8'd139, 8'd63, 8'd129, 8'd141, 8'd136, 8'd149, 8'd87, 8'd93, 8'd135, 8'd103, 8'd147, 8'd150, 8'd57, 8'd140, 8'd105, 8'd130, 8'd100, 8'd90, 8'd107, 8'd86, 8'd119, 8'd104, 8'd78, 8'd112, 8'd114, 8'd119, 8'd152, 8'd115, 8'd128, 8'd85, 8'd147, 8'd99, 8'd131, 8'd133, 8'd143, 8'd164, 8'd96, 8'd168, 8'd110, 8'd125, 8'd90, 8'd77, 8'd98, 8'd138, 8'd141, 8'd120, 8'd89, 8'd91, 8'd107, 8'd145, 8'd166, 8'd114, 8'd76, 8'd114, 8'd95, 8'd155, 8'd78, 8'd73, 8'd127, 8'd136, 8'd166, 8'd85, 8'd169, 8'd107, 8'd146, 8'd100, 8'd81, 8'd78, 8'd126, 8'd94, 8'd122, 8'd106, 8'd101, 8'd88, 8'd83, 8'd132, 8'd72, 8'd63, 8'd72, 8'd146, 8'd90, 8'd72, 8'd69, 8'd68, 8'd126, 8'd86, 8'd79, 8'd80, 8'd107, 8'd78, 8'd80, 8'd91, 8'd93, 8'd166, 8'd129, 8'd144, 8'd116, 8'd126, 8'd75, 8'd116, 8'd161, 8'd110, 8'd139, 8'd146, 8'd76, 8'd131, 8'd70, 8'd88, 8'd133, 8'd98, 8'd112, 8'd111, 8'd152, 8'd148, 8'd82, 8'd121, 8'd159, 8'd162, 8'd118, 8'd142, 8'd94, 8'd127, 8'd167, 8'd79, 8'd74, 8'd109, 8'd81, 8'd98, 8'd75, 8'd166, 8'd102, 8'd108, 8'd103, 8'd116, 8'd112, 8'd108, 8'd126, 8'd158, 8'd86, 8'd79, 8'd141, 8'd108, 8'd79, 8'd132, 8'd157, 8'd113})
) cell_0_62 (
    .clk(clk),
    .input_index(index_0_61_62),
    .input_value(value_0_61_62),
    .input_result(result_0_61_62),
    .input_enable(enable_0_61_62),
    .output_index(index_0_62_63),
    .output_value(value_0_62_63),
    .output_result(result_0_62_63),
    .output_enable(enable_0_62_63)
);

wire [10-1:0] index_0_63_64;
wire [`DATA_WIDTH-1:0] value_0_63_64;
wire [`DATA_WIDTH*4:0] result_0_63_64;
wire enable_0_63_64;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd117, 8'd145, 8'd168, 8'd99, 8'd128, 8'd72, 8'd69, 8'd154, 8'd148, 8'd135, 8'd110, 8'd129, 8'd133, 8'd154, 8'd128, 8'd166, 8'd139, 8'd84, 8'd145, 8'd106, 8'd82, 8'd123, 8'd133, 8'd106, 8'd116, 8'd149, 8'd152, 8'd164, 8'd149, 8'd137, 8'd88, 8'd116, 8'd156, 8'd164, 8'd129, 8'd111, 8'd118, 8'd138, 8'd175, 8'd117, 8'd130, 8'd124, 8'd173, 8'd159, 8'd128, 8'd123, 8'd147, 8'd192, 8'd181, 8'd161, 8'd121, 8'd141, 8'd104, 8'd126, 8'd130, 8'd160, 8'd74, 8'd127, 8'd68, 8'd70, 8'd149, 8'd99, 8'd150, 8'd130, 8'd165, 8'd129, 8'd100, 8'd84, 8'd124, 8'd125, 8'd95, 8'd137, 8'd161, 8'd122, 8'd76, 8'd169, 8'd111, 8'd127, 8'd159, 8'd123, 8'd113, 8'd159, 8'd142, 8'd138, 8'd151, 8'd155, 8'd97, 8'd127, 8'd101, 8'd79, 8'd175, 8'd133, 8'd95, 8'd87, 8'd134, 8'd103, 8'd119, 8'd145, 8'd165, 8'd96, 8'd91, 8'd175, 8'd77, 8'd109, 8'd143, 8'd90, 8'd127, 8'd133, 8'd137, 8'd97, 8'd152, 8'd83, 8'd143, 8'd104, 8'd86, 8'd147, 8'd124, 8'd146, 8'd165, 8'd116, 8'd105, 8'd82, 8'd82, 8'd118, 8'd115, 8'd87, 8'd146, 8'd162, 8'd93, 8'd169, 8'd121, 8'd130, 8'd104, 8'd84, 8'd138, 8'd98, 8'd113, 8'd70, 8'd79, 8'd159, 8'd108, 8'd140, 8'd162, 8'd122, 8'd141, 8'd159, 8'd133, 8'd107, 8'd101, 8'd152, 8'd166, 8'd140, 8'd142, 8'd108, 8'd123, 8'd140, 8'd145, 8'd156, 8'd122, 8'd118, 8'd90, 8'd87, 8'd168, 8'd72, 8'd82, 8'd149, 8'd123, 8'd75, 8'd124, 8'd56, 8'd79, 8'd148, 8'd65, 8'd96, 8'd140, 8'd89, 8'd129, 8'd78, 8'd72, 8'd89, 8'd84, 8'd126, 8'd134, 8'd68, 8'd112, 8'd124, 8'd85, 8'd107, 8'd143, 8'd126, 8'd125, 8'd120, 8'd73, 8'd67, 8'd140, 8'd89, 8'd125, 8'd114, 8'd115, 8'd85, 8'd99, 8'd150, 8'd150, 8'd158, 8'd147, 8'd85, 8'd120, 8'd156, 8'd112, 8'd117, 8'd119, 8'd92, 8'd104, 8'd143, 8'd75, 8'd161, 8'd170, 8'd170, 8'd70, 8'd73, 8'd80, 8'd108, 8'd67, 8'd81, 8'd111, 8'd74, 8'd99, 8'd114, 8'd144, 8'd157, 8'd94, 8'd127, 8'd90, 8'd105, 8'd82, 8'd153, 8'd153, 8'd150, 8'd98, 8'd101, 8'd61, 8'd115, 8'd157, 8'd74, 8'd89, 8'd142, 8'd92, 8'd65, 8'd130, 8'd85, 8'd75, 8'd174, 8'd111, 8'd128, 8'd57, 8'd48, 8'd72, 8'd152, 8'd70, 8'd134, 8'd119, 8'd83, 8'd60, 8'd114, 8'd114, 8'd149, 8'd142, 8'd107, 8'd148, 8'd147, 8'd148, 8'd121, 8'd83, 8'd121, 8'd59, 8'd151, 8'd150, 8'd154, 8'd115, 8'd141, 8'd105, 8'd158, 8'd50, 8'd60, 8'd67, 8'd142, 8'd72, 8'd77, 8'd106, 8'd135, 8'd135, 8'd111, 8'd152, 8'd79, 8'd83, 8'd104, 8'd83, 8'd132, 8'd140, 8'd134, 8'd93, 8'd147, 8'd135, 8'd112, 8'd158, 8'd76, 8'd145, 8'd141, 8'd90, 8'd130, 8'd148, 8'd108, 8'd89, 8'd114, 8'd93, 8'd68, 8'd54, 8'd112, 8'd156, 8'd95, 8'd113, 8'd87, 8'd137, 8'd119, 8'd118, 8'd143, 8'd100, 8'd145, 8'd94, 8'd141, 8'd92, 8'd94, 8'd83, 8'd150, 8'd151, 8'd84, 8'd140, 8'd84, 8'd97, 8'd138, 8'd62, 8'd74, 8'd125, 8'd136, 8'd131, 8'd127, 8'd105, 8'd111, 8'd129, 8'd115, 8'd103, 8'd134, 8'd64, 8'd83, 8'd73, 8'd109, 8'd106, 8'd86, 8'd142, 8'd150, 8'd135, 8'd61, 8'd125, 8'd159, 8'd80, 8'd171, 8'd156, 8'd102, 8'd67, 8'd124, 8'd117, 8'd116, 8'd129, 8'd117, 8'd118, 8'd147, 8'd107, 8'd105, 8'd186, 8'd149, 8'd109, 8'd80, 8'd137, 8'd118, 8'd145, 8'd147, 8'd110, 8'd98, 8'd166, 8'd58, 8'd151, 8'd127, 8'd119, 8'd140, 8'd145, 8'd115, 8'd162, 8'd131, 8'd124, 8'd94, 8'd113, 8'd162, 8'd93, 8'd154, 8'd116, 8'd112, 8'd109, 8'd125, 8'd92, 8'd57, 8'd102, 8'd81, 8'd62, 8'd101, 8'd127, 8'd89, 8'd142, 8'd100, 8'd151, 8'd150, 8'd154, 8'd89, 8'd79, 8'd94, 8'd120, 8'd194, 8'd135, 8'd118, 8'd96, 8'd159, 8'd162, 8'd146, 8'd149, 8'd204, 8'd170, 8'd120, 8'd98, 8'd86, 8'd86, 8'd81, 8'd152, 8'd93, 8'd131, 8'd148, 8'd134, 8'd72, 8'd158, 8'd105, 8'd111, 8'd76, 8'd93, 8'd128, 8'd128, 8'd130, 8'd118, 8'd98, 8'd104, 8'd137, 8'd102, 8'd172, 8'd154, 8'd105, 8'd106, 8'd140, 8'd106, 8'd122, 8'd80, 8'd92, 8'd165, 8'd132, 8'd146, 8'd120, 8'd119, 8'd109, 8'd141, 8'd92, 8'd169, 8'd95, 8'd84, 8'd74, 8'd121, 8'd118, 8'd145, 8'd138, 8'd111, 8'd131, 8'd108, 8'd84, 8'd170, 8'd116, 8'd90, 8'd91, 8'd163, 8'd116, 8'd138, 8'd105, 8'd93, 8'd145, 8'd132, 8'd159, 8'd154, 8'd73, 8'd68, 8'd82, 8'd106, 8'd103, 8'd85, 8'd47, 8'd85, 8'd107, 8'd103, 8'd178, 8'd156, 8'd185, 8'd154, 8'd133, 8'd127, 8'd100, 8'd98, 8'd94, 8'd140, 8'd96, 8'd93, 8'd94, 8'd152, 8'd144, 8'd179, 8'd128, 8'd85, 8'd108, 8'd124, 8'd107, 8'd147, 8'd146, 8'd68, 8'd99, 8'd121, 8'd162, 8'd88, 8'd104, 8'd84, 8'd167, 8'd132, 8'd90, 8'd154, 8'd114, 8'd144, 8'd138, 8'd137, 8'd106, 8'd143, 8'd144, 8'd129, 8'd152, 8'd125, 8'd123, 8'd72, 8'd67, 8'd80, 8'd161, 8'd130, 8'd79, 8'd87, 8'd73, 8'd84, 8'd132, 8'd139, 8'd119, 8'd125, 8'd157, 8'd107, 8'd98, 8'd144, 8'd183, 8'd137, 8'd103, 8'd87, 8'd125, 8'd101, 8'd115, 8'd84, 8'd136, 8'd73, 8'd112, 8'd138, 8'd83, 8'd75, 8'd83, 8'd77, 8'd149, 8'd60, 8'd114, 8'd142, 8'd78, 8'd69, 8'd79, 8'd108, 8'd168, 8'd142, 8'd157, 8'd130, 8'd112, 8'd156, 8'd128, 8'd123, 8'd85, 8'd150, 8'd117, 8'd81, 8'd65, 8'd66, 8'd67, 8'd109, 8'd131, 8'd106, 8'd70, 8'd126, 8'd64, 8'd102, 8'd116, 8'd48, 8'd133, 8'd89, 8'd134, 8'd123, 8'd109, 8'd155, 8'd129, 8'd93, 8'd121, 8'd132, 8'd125, 8'd126, 8'd114, 8'd97, 8'd56, 8'd157, 8'd138, 8'd99, 8'd132, 8'd104, 8'd130, 8'd112, 8'd136, 8'd130, 8'd116, 8'd108, 8'd71, 8'd76, 8'd137, 8'd141, 8'd117, 8'd109, 8'd144, 8'd117, 8'd98, 8'd156, 8'd166, 8'd137, 8'd155, 8'd155, 8'd100, 8'd112, 8'd134, 8'd91, 8'd123, 8'd91, 8'd74, 8'd127, 8'd158, 8'd92, 8'd169, 8'd74, 8'd117, 8'd158, 8'd161, 8'd83, 8'd100, 8'd93, 8'd102, 8'd84, 8'd124, 8'd80, 8'd83, 8'd78, 8'd74, 8'd83, 8'd58, 8'd68, 8'd113, 8'd97, 8'd68, 8'd101, 8'd147, 8'd151, 8'd148, 8'd111, 8'd113, 8'd126, 8'd89, 8'd153, 8'd160, 8'd114, 8'd77, 8'd86, 8'd75, 8'd139, 8'd129, 8'd127, 8'd123, 8'd76, 8'd148, 8'd99, 8'd163, 8'd147, 8'd98, 8'd83, 8'd112, 8'd97, 8'd93, 8'd141, 8'd84, 8'd164, 8'd96, 8'd86, 8'd73, 8'd112, 8'd130, 8'd96, 8'd111, 8'd70, 8'd77, 8'd119, 8'd147, 8'd118, 8'd107, 8'd145, 8'd89, 8'd127, 8'd152, 8'd158, 8'd168, 8'd91, 8'd140, 8'd165, 8'd106, 8'd160, 8'd106, 8'd88, 8'd86, 8'd89, 8'd153, 8'd79, 8'd103, 8'd84, 8'd138, 8'd151, 8'd122, 8'd95, 8'd144, 8'd122, 8'd167, 8'd154, 8'd168, 8'd115, 8'd118, 8'd121, 8'd135, 8'd76, 8'd86, 8'd126, 8'd95, 8'd92, 8'd97, 8'd138, 8'd103, 8'd117, 8'd127, 8'd169, 8'd88, 8'd107, 8'd95, 8'd107, 8'd130})
) cell_0_63 (
    .clk(clk),
    .input_index(index_0_62_63),
    .input_value(value_0_62_63),
    .input_result(result_0_62_63),
    .input_enable(enable_0_62_63),
    .output_index(index_0_63_64),
    .output_value(value_0_63_64),
    .output_result(result_0_63_64),
    .output_enable(enable_0_63_64)
);

wire [10-1:0] index_0_64_65;
wire [`DATA_WIDTH-1:0] value_0_64_65;
wire [`DATA_WIDTH*4:0] result_0_64_65;
wire enable_0_64_65;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd136, 8'd105, 8'd74, 8'd117, 8'd110, 8'd81, 8'd147, 8'd134, 8'd112, 8'd67, 8'd65, 8'd117, 8'd96, 8'd122, 8'd124, 8'd109, 8'd130, 8'd121, 8'd84, 8'd121, 8'd130, 8'd137, 8'd108, 8'd130, 8'd166, 8'd109, 8'd106, 8'd141, 8'd88, 8'd90, 8'd167, 8'd96, 8'd123, 8'd107, 8'd90, 8'd65, 8'd129, 8'd37, 8'd50, 8'd38, 8'd76, 8'd64, 8'd38, 8'd115, 8'd80, 8'd62, 8'd81, 8'd102, 8'd91, 8'd171, 8'd116, 8'd140, 8'd172, 8'd85, 8'd73, 8'd145, 8'd114, 8'd136, 8'd115, 8'd148, 8'd87, 8'd52, 8'd66, 8'd86, 8'd51, 8'd65, 8'd46, 8'd134, 8'd101, 8'd148, 8'd95, 8'd149, 8'd112, 8'd122, 8'd84, 8'd156, 8'd114, 8'd124, 8'd143, 8'd167, 8'd160, 8'd157, 8'd94, 8'd162, 8'd117, 8'd134, 8'd121, 8'd120, 8'd156, 8'd135, 8'd129, 8'd129, 8'd126, 8'd153, 8'd82, 8'd69, 8'd74, 8'd69, 8'd128, 8'd102, 8'd74, 8'd162, 8'd104, 8'd132, 8'd100, 8'd102, 8'd169, 8'd164, 8'd134, 8'd126, 8'd71, 8'd78, 8'd73, 8'd128, 8'd129, 8'd105, 8'd154, 8'd121, 8'd115, 8'd163, 8'd156, 8'd101, 8'd82, 8'd62, 8'd52, 8'd106, 8'd117, 8'd86, 8'd68, 8'd66, 8'd144, 8'd139, 8'd80, 8'd130, 8'd74, 8'd177, 8'd86, 8'd101, 8'd78, 8'd143, 8'd131, 8'd137, 8'd83, 8'd138, 8'd156, 8'd102, 8'd174, 8'd117, 8'd153, 8'd88, 8'd92, 8'd85, 8'd77, 8'd93, 8'd138, 8'd72, 8'd72, 8'd134, 8'd124, 8'd159, 8'd121, 8'd134, 8'd150, 8'd155, 8'd170, 8'd133, 8'd88, 8'd88, 8'd134, 8'd81, 8'd158, 8'd127, 8'd113, 8'd119, 8'd73, 8'd168, 8'd183, 8'd128, 8'd116, 8'd133, 8'd135, 8'd178, 8'd108, 8'd181, 8'd147, 8'd116, 8'd168, 8'd68, 8'd55, 8'd75, 8'd83, 8'd81, 8'd91, 8'd94, 8'd81, 8'd135, 8'd108, 8'd95, 8'd193, 8'd107, 8'd119, 8'd78, 8'd166, 8'd155, 8'd144, 8'd190, 8'd183, 8'd186, 8'd154, 8'd152, 8'd153, 8'd169, 8'd166, 8'd100, 8'd175, 8'd110, 8'd129, 8'd88, 8'd61, 8'd171, 8'd103, 8'd79, 8'd92, 8'd82, 8'd104, 8'd94, 8'd167, 8'd138, 8'd185, 8'd133, 8'd182, 8'd188, 8'd184, 8'd186, 8'd140, 8'd165, 8'd142, 8'd177, 8'd162, 8'd132, 8'd125, 8'd101, 8'd108, 8'd154, 8'd103, 8'd135, 8'd131, 8'd98, 8'd147, 8'd139, 8'd125, 8'd121, 8'd93, 8'd147, 8'd194, 8'd186, 8'd193, 8'd92, 8'd188, 8'd112, 8'd123, 8'd104, 8'd182, 8'd165, 8'd89, 8'd114, 8'd167, 8'd152, 8'd192, 8'd166, 8'd127, 8'd176, 8'd174, 8'd109, 8'd132, 8'd113, 8'd175, 8'd88, 8'd160, 8'd143, 8'd77, 8'd179, 8'd140, 8'd172, 8'd140, 8'd159, 8'd92, 8'd109, 8'd130, 8'd161, 8'd122, 8'd122, 8'd124, 8'd99, 8'd144, 8'd104, 8'd117, 8'd183, 8'd121, 8'd161, 8'd146, 8'd124, 8'd87, 8'd136, 8'd118, 8'd97, 8'd119, 8'd132, 8'd109, 8'd167, 8'd218, 8'd178, 8'd102, 8'd89, 8'd167, 8'd129, 8'd167, 8'd124, 8'd144, 8'd115, 8'd105, 8'd85, 8'd96, 8'd138, 8'd187, 8'd195, 8'd91, 8'd109, 8'd191, 8'd100, 8'd139, 8'd131, 8'd92, 8'd164, 8'd62, 8'd122, 8'd138, 8'd157, 8'd167, 8'd145, 8'd133, 8'd147, 8'd136, 8'd110, 8'd122, 8'd94, 8'd125, 8'd206, 8'd173, 8'd103, 8'd112, 8'd135, 8'd210, 8'd162, 8'd178, 8'd153, 8'd152, 8'd188, 8'd168, 8'd114, 8'd157, 8'd83, 8'd95, 8'd153, 8'd166, 8'd144, 8'd153, 8'd154, 8'd103, 8'd184, 8'd122, 8'd163, 8'd163, 8'd141, 8'd159, 8'd125, 8'd130, 8'd127, 8'd94, 8'd185, 8'd123, 8'd144, 8'd171, 8'd99, 8'd113, 8'd163, 8'd72, 8'd71, 8'd105, 8'd101, 8'd136, 8'd107, 8'd105, 8'd117, 8'd128, 8'd216, 8'd157, 8'd161, 8'd144, 8'd129, 8'd143, 8'd121, 8'd122, 8'd121, 8'd91, 8'd95, 8'd142, 8'd116, 8'd176, 8'd131, 8'd136, 8'd109, 8'd126, 8'd67, 8'd109, 8'd125, 8'd68, 8'd106, 8'd62, 8'd114, 8'd139, 8'd146, 8'd96, 8'd115, 8'd110, 8'd154, 8'd116, 8'd132, 8'd126, 8'd133, 8'd102, 8'd172, 8'd126, 8'd99, 8'd139, 8'd93, 8'd68, 8'd92, 8'd93, 8'd62, 8'd66, 8'd114, 8'd135, 8'd110, 8'd116, 8'd67, 8'd152, 8'd102, 8'd78, 8'd63, 8'd52, 8'd97, 8'd134, 8'd119, 8'd95, 8'd156, 8'd81, 8'd67, 8'd77, 8'd67, 8'd94, 8'd69, 8'd69, 8'd96, 8'd97, 8'd63, 8'd105, 8'd113, 8'd42, 8'd57, 8'd104, 8'd125, 8'd158, 8'd141, 8'd70, 8'd96, 8'd89, 8'd102, 8'd33, 8'd54, 8'd108, 8'd110, 8'd105, 8'd144, 8'd70, 8'd55, 8'd66, 8'd81, 8'd83, 8'd91, 8'd52, 8'd79, 8'd117, 8'd143, 8'd96, 8'd67, 8'd140, 8'd147, 8'd148, 8'd71, 8'd114, 8'd140, 8'd64, 8'd96, 8'd111, 8'd83, 8'd84, 8'd30, 8'd96, 8'd82, 8'd95, 8'd85, 8'd40, 8'd88, 8'd104, 8'd107, 8'd123, 8'd111, 8'd124, 8'd129, 8'd149, 8'd127, 8'd169, 8'd76, 8'd166, 8'd158, 8'd79, 8'd176, 8'd148, 8'd122, 8'd145, 8'd106, 8'd56, 8'd93, 8'd45, 8'd6, 8'd49, 8'd71, 8'd88, 8'd60, 8'd84, 8'd69, 8'd100, 8'd117, 8'd113, 8'd88, 8'd110, 8'd166, 8'd143, 8'd178, 8'd142, 8'd167, 8'd88, 8'd78, 8'd163, 8'd118, 8'd133, 8'd117, 8'd138, 8'd93, 8'd117, 8'd104, 8'd54, 8'd84, 8'd27, 8'd73, 8'd78, 8'd46, 8'd105, 8'd75, 8'd128, 8'd163, 8'd176, 8'd123, 8'd134, 8'd131, 8'd94, 8'd175, 8'd158, 8'd113, 8'd179, 8'd124, 8'd170, 8'd158, 8'd80, 8'd174, 8'd91, 8'd89, 8'd155, 8'd80, 8'd117, 8'd130, 8'd48, 8'd137, 8'd71, 8'd84, 8'd92, 8'd146, 8'd163, 8'd103, 8'd178, 8'd151, 8'd160, 8'd109, 8'd117, 8'd113, 8'd123, 8'd144, 8'd142, 8'd181, 8'd148, 8'd174, 8'd102, 8'd87, 8'd126, 8'd95, 8'd167, 8'd105, 8'd109, 8'd153, 8'd120, 8'd146, 8'd104, 8'd159, 8'd84, 8'd135, 8'd130, 8'd155, 8'd88, 8'd94, 8'd95, 8'd134, 8'd168, 8'd170, 8'd168, 8'd132, 8'd177, 8'd93, 8'd109, 8'd179, 8'd94, 8'd155, 8'd78, 8'd125, 8'd110, 8'd142, 8'd88, 8'd137, 8'd138, 8'd91, 8'd94, 8'd121, 8'd188, 8'd100, 8'd158, 8'd91, 8'd101, 8'd110, 8'd155, 8'd100, 8'd145, 8'd172, 8'd133, 8'd131, 8'd153, 8'd168, 8'd120, 8'd93, 8'd141, 8'd140, 8'd81, 8'd113, 8'd101, 8'd109, 8'd149, 8'd186, 8'd152, 8'd145, 8'd115, 8'd163, 8'd123, 8'd204, 8'd114, 8'd149, 8'd124, 8'd176, 8'd197, 8'd153, 8'd156, 8'd128, 8'd204, 8'd133, 8'd149, 8'd158, 8'd166, 8'd78, 8'd80, 8'd81, 8'd131, 8'd166, 8'd131, 8'd114, 8'd155, 8'd113, 8'd133, 8'd176, 8'd200, 8'd149, 8'd158, 8'd192, 8'd177, 8'd189, 8'd169, 8'd124, 8'd134, 8'd213, 8'd162, 8'd195, 8'd147, 8'd207, 8'd112, 8'd116, 8'd105, 8'd99, 8'd149, 8'd133, 8'd156, 8'd140, 8'd100, 8'd142, 8'd89, 8'd147, 8'd108, 8'd107, 8'd121, 8'd97, 8'd155, 8'd97, 8'd178, 8'd133, 8'd95, 8'd140, 8'd178, 8'd151, 8'd154, 8'd98, 8'd129, 8'd171, 8'd112, 8'd163, 8'd90, 8'd137, 8'd102, 8'd74, 8'd87, 8'd117, 8'd89, 8'd119, 8'd73, 8'd107, 8'd99, 8'd168, 8'd143, 8'd70, 8'd134, 8'd133, 8'd79, 8'd167, 8'd158, 8'd129, 8'd88, 8'd105, 8'd106, 8'd133, 8'd132, 8'd96, 8'd83, 8'd138, 8'd164, 8'd83, 8'd87, 8'd102, 8'd161, 8'd159})
) cell_0_64 (
    .clk(clk),
    .input_index(index_0_63_64),
    .input_value(value_0_63_64),
    .input_result(result_0_63_64),
    .input_enable(enable_0_63_64),
    .output_index(index_0_64_65),
    .output_value(value_0_64_65),
    .output_result(result_0_64_65),
    .output_enable(enable_0_64_65)
);

wire [10-1:0] index_0_65_66;
wire [`DATA_WIDTH-1:0] value_0_65_66;
wire [`DATA_WIDTH*4:0] result_0_65_66;
wire enable_0_65_66;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd134, 8'd116, 8'd90, 8'd112, 8'd136, 8'd114, 8'd90, 8'd168, 8'd115, 8'd75, 8'd98, 8'd88, 8'd78, 8'd105, 8'd125, 8'd105, 8'd130, 8'd61, 8'd89, 8'd90, 8'd95, 8'd111, 8'd140, 8'd166, 8'd160, 8'd77, 8'd153, 8'd96, 8'd145, 8'd83, 8'd117, 8'd99, 8'd93, 8'd136, 8'd107, 8'd169, 8'd103, 8'd76, 8'd73, 8'd77, 8'd147, 8'd117, 8'd90, 8'd173, 8'd93, 8'd92, 8'd174, 8'd179, 8'd143, 8'd145, 8'd122, 8'd175, 8'd134, 8'd134, 8'd101, 8'd93, 8'd125, 8'd119, 8'd87, 8'd128, 8'd110, 8'd152, 8'd120, 8'd184, 8'd98, 8'd130, 8'd175, 8'd151, 8'd89, 8'd94, 8'd170, 8'd133, 8'd189, 8'd134, 8'd137, 8'd198, 8'd166, 8'd177, 8'd156, 8'd158, 8'd156, 8'd148, 8'd83, 8'd84, 8'd93, 8'd113, 8'd144, 8'd155, 8'd127, 8'd178, 8'd192, 8'd173, 8'd128, 8'd97, 8'd94, 8'd114, 8'd144, 8'd65, 8'd90, 8'd115, 8'd104, 8'd95, 8'd169, 8'd175, 8'd171, 8'd142, 8'd133, 8'd116, 8'd169, 8'd136, 8'd73, 8'd84, 8'd149, 8'd157, 8'd119, 8'd135, 8'd132, 8'd164, 8'd167, 8'd112, 8'd115, 8'd123, 8'd116, 8'd61, 8'd147, 8'd97, 8'd47, 8'd92, 8'd118, 8'd92, 8'd142, 8'd128, 8'd155, 8'd95, 8'd152, 8'd177, 8'd158, 8'd122, 8'd133, 8'd121, 8'd135, 8'd154, 8'd136, 8'd164, 8'd100, 8'd153, 8'd91, 8'd139, 8'd170, 8'd123, 8'd132, 8'd159, 8'd140, 8'd116, 8'd129, 8'd151, 8'd157, 8'd64, 8'd80, 8'd84, 8'd60, 8'd67, 8'd84, 8'd164, 8'd105, 8'd149, 8'd146, 8'd85, 8'd132, 8'd105, 8'd126, 8'd181, 8'd91, 8'd82, 8'd74, 8'd95, 8'd82, 8'd134, 8'd89, 8'd168, 8'd103, 8'd87, 8'd87, 8'd84, 8'd119, 8'd128, 8'd96, 8'd96, 8'd72, 8'd128, 8'd118, 8'd118, 8'd148, 8'd158, 8'd117, 8'd105, 8'd89, 8'd169, 8'd159, 8'd95, 8'd117, 8'd79, 8'd136, 8'd156, 8'd144, 8'd77, 8'd86, 8'd124, 8'd124, 8'd123, 8'd71, 8'd150, 8'd139, 8'd114, 8'd75, 8'd57, 8'd145, 8'd129, 8'd125, 8'd135, 8'd103, 8'd158, 8'd141, 8'd82, 8'd172, 8'd141, 8'd170, 8'd139, 8'd64, 8'd87, 8'd129, 8'd169, 8'd132, 8'd126, 8'd168, 8'd160, 8'd104, 8'd133, 8'd134, 8'd79, 8'd86, 8'd111, 8'd80, 8'd136, 8'd114, 8'd96, 8'd82, 8'd157, 8'd171, 8'd132, 8'd83, 8'd90, 8'd92, 8'd142, 8'd78, 8'd140, 8'd157, 8'd103, 8'd142, 8'd170, 8'd94, 8'd106, 8'd125, 8'd91, 8'd144, 8'd91, 8'd136, 8'd127, 8'd134, 8'd93, 8'd56, 8'd55, 8'd160, 8'd119, 8'd110, 8'd147, 8'd118, 8'd124, 8'd83, 8'd111, 8'd69, 8'd174, 8'd89, 8'd69, 8'd80, 8'd149, 8'd109, 8'd94, 8'd156, 8'd132, 8'd133, 8'd148, 8'd179, 8'd141, 8'd101, 8'd62, 8'd97, 8'd69, 8'd125, 8'd145, 8'd149, 8'd78, 8'd162, 8'd152, 8'd105, 8'd105, 8'd122, 8'd156, 8'd143, 8'd109, 8'd143, 8'd63, 8'd70, 8'd144, 8'd92, 8'd139, 8'd140, 8'd130, 8'd142, 8'd144, 8'd152, 8'd153, 8'd140, 8'd140, 8'd168, 8'd122, 8'd84, 8'd118, 8'd111, 8'd106, 8'd157, 8'd149, 8'd76, 8'd148, 8'd74, 8'd82, 8'd124, 8'd137, 8'd142, 8'd62, 8'd97, 8'd94, 8'd94, 8'd116, 8'd82, 8'd107, 8'd129, 8'd189, 8'd139, 8'd70, 8'd110, 8'd94, 8'd173, 8'd99, 8'd87, 8'd125, 8'd157, 8'd140, 8'd110, 8'd164, 8'd107, 8'd71, 8'd81, 8'd134, 8'd121, 8'd72, 8'd120, 8'd95, 8'd82, 8'd131, 8'd120, 8'd181, 8'd132, 8'd102, 8'd152, 8'd167, 8'd130, 8'd85, 8'd96, 8'd156, 8'd145, 8'd181, 8'd121, 8'd146, 8'd103, 8'd126, 8'd90, 8'd135, 8'd156, 8'd61, 8'd150, 8'd168, 8'd111, 8'd143, 8'd61, 8'd65, 8'd41, 8'd87, 8'd161, 8'd101, 8'd178, 8'd180, 8'd186, 8'd140, 8'd88, 8'd169, 8'd135, 8'd165, 8'd186, 8'd146, 8'd122, 8'd161, 8'd164, 8'd104, 8'd126, 8'd158, 8'd111, 8'd47, 8'd132, 8'd147, 8'd119, 8'd120, 8'd127, 8'd17, 8'd69, 8'd93, 8'd68, 8'd139, 8'd140, 8'd155, 8'd165, 8'd147, 8'd170, 8'd141, 8'd104, 8'd139, 8'd130, 8'd106, 8'd92, 8'd152, 8'd101, 8'd133, 8'd113, 8'd156, 8'd141, 8'd49, 8'd52, 8'd88, 8'd157, 8'd141, 8'd161, 8'd62, 8'd100, 8'd102, 8'd104, 8'd89, 8'd76, 8'd79, 8'd156, 8'd99, 8'd95, 8'd61, 8'd154, 8'd135, 8'd128, 8'd151, 8'd140, 8'd150, 8'd157, 8'd156, 8'd160, 8'd121, 8'd90, 8'd81, 8'd117, 8'd161, 8'd121, 8'd99, 8'd127, 8'd90, 8'd67, 8'd66, 8'd131, 8'd121, 8'd125, 8'd101, 8'd113, 8'd143, 8'd77, 8'd95, 8'd65, 8'd108, 8'd124, 8'd141, 8'd113, 8'd93, 8'd98, 8'd158, 8'd69, 8'd47, 8'd65, 8'd66, 8'd137, 8'd118, 8'd117, 8'd121, 8'd124, 8'd133, 8'd144, 8'd114, 8'd73, 8'd74, 8'd88, 8'd134, 8'd125, 8'd137, 8'd157, 8'd97, 8'd138, 8'd84, 8'd126, 8'd142, 8'd94, 8'd110, 8'd104, 8'd76, 8'd119, 8'd73, 8'd81, 8'd123, 8'd94, 8'd86, 8'd71, 8'd165, 8'd180, 8'd92, 8'd144, 8'd76, 8'd77, 8'd114, 8'd105, 8'd70, 8'd116, 8'd115, 8'd164, 8'd89, 8'd162, 8'd133, 8'd88, 8'd147, 8'd125, 8'd159, 8'd64, 8'd143, 8'd145, 8'd49, 8'd80, 8'd131, 8'd129, 8'd126, 8'd113, 8'd84, 8'd173, 8'd135, 8'd98, 8'd114, 8'd107, 8'd110, 8'd126, 8'd149, 8'd82, 8'd172, 8'd127, 8'd128, 8'd150, 8'd117, 8'd172, 8'd155, 8'd120, 8'd91, 8'd138, 8'd98, 8'd110, 8'd113, 8'd135, 8'd98, 8'd94, 8'd161, 8'd177, 8'd152, 8'd113, 8'd179, 8'd157, 8'd78, 8'd117, 8'd149, 8'd132, 8'd114, 8'd144, 8'd152, 8'd96, 8'd116, 8'd166, 8'd118, 8'd120, 8'd109, 8'd149, 8'd116, 8'd160, 8'd134, 8'd92, 8'd142, 8'd79, 8'd82, 8'd148, 8'd130, 8'd91, 8'd175, 8'd111, 8'd91, 8'd93, 8'd156, 8'd122, 8'd151, 8'd93, 8'd153, 8'd95, 8'd72, 8'd113, 8'd136, 8'd70, 8'd65, 8'd123, 8'd148, 8'd149, 8'd153, 8'd93, 8'd90, 8'd120, 8'd151, 8'd123, 8'd116, 8'd153, 8'd73, 8'd169, 8'd129, 8'd167, 8'd168, 8'd88, 8'd123, 8'd135, 8'd90, 8'd128, 8'd82, 8'd118, 8'd129, 8'd50, 8'd143, 8'd109, 8'd139, 8'd140, 8'd70, 8'd153, 8'd94, 8'd130, 8'd146, 8'd128, 8'd80, 8'd88, 8'd85, 8'd118, 8'd151, 8'd159, 8'd93, 8'd160, 8'd89, 8'd112, 8'd142, 8'd97, 8'd111, 8'd104, 8'd126, 8'd102, 8'd119, 8'd72, 8'd83, 8'd67, 8'd120, 8'd78, 8'd101, 8'd158, 8'd151, 8'd138, 8'd66, 8'd101, 8'd169, 8'd151, 8'd146, 8'd164, 8'd115, 8'd138, 8'd144, 8'd153, 8'd136, 8'd93, 8'd139, 8'd154, 8'd99, 8'd125, 8'd152, 8'd141, 8'd101, 8'd88, 8'd138, 8'd82, 8'd84, 8'd82, 8'd38, 8'd145, 8'd100, 8'd83, 8'd76, 8'd98, 8'd78, 8'd110, 8'd154, 8'd107, 8'd143, 8'd87, 8'd141, 8'd161, 8'd113, 8'd151, 8'd116, 8'd120, 8'd116, 8'd63, 8'd113, 8'd74, 8'd131, 8'd63, 8'd100, 8'd120, 8'd124, 8'd89, 8'd140, 8'd125, 8'd118, 8'd102, 8'd63, 8'd123, 8'd114, 8'd117, 8'd83, 8'd104, 8'd143, 8'd123, 8'd96, 8'd131, 8'd129, 8'd98, 8'd161, 8'd134, 8'd133, 8'd105, 8'd103, 8'd167, 8'd79, 8'd97, 8'd132, 8'd142, 8'd93, 8'd86, 8'd103, 8'd79, 8'd160, 8'd160, 8'd109, 8'd124, 8'd129, 8'd118, 8'd117, 8'd162, 8'd128})
) cell_0_65 (
    .clk(clk),
    .input_index(index_0_64_65),
    .input_value(value_0_64_65),
    .input_result(result_0_64_65),
    .input_enable(enable_0_64_65),
    .output_index(index_0_65_66),
    .output_value(value_0_65_66),
    .output_result(result_0_65_66),
    .output_enable(enable_0_65_66)
);

wire [10-1:0] index_0_66_67;
wire [`DATA_WIDTH-1:0] value_0_66_67;
wire [`DATA_WIDTH*4:0] result_0_66_67;
wire enable_0_66_67;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd165, 8'd98, 8'd75, 8'd132, 8'd137, 8'd154, 8'd123, 8'd111, 8'd143, 8'd148, 8'd74, 8'd120, 8'd111, 8'd104, 8'd103, 8'd78, 8'd97, 8'd84, 8'd123, 8'd93, 8'd145, 8'd98, 8'd121, 8'd122, 8'd71, 8'd170, 8'd136, 8'd111, 8'd170, 8'd114, 8'd69, 8'd87, 8'd121, 8'd147, 8'd171, 8'd125, 8'd99, 8'd127, 8'd125, 8'd98, 8'd161, 8'd140, 8'd169, 8'd187, 8'd125, 8'd169, 8'd160, 8'd185, 8'd166, 8'd109, 8'd185, 8'd146, 8'd147, 8'd139, 8'd82, 8'd151, 8'd101, 8'd135, 8'd139, 8'd184, 8'd91, 8'd92, 8'd113, 8'd177, 8'd125, 8'd145, 8'd113, 8'd114, 8'd187, 8'd126, 8'd123, 8'd131, 8'd108, 8'd182, 8'd101, 8'd102, 8'd175, 8'd107, 8'd150, 8'd86, 8'd131, 8'd105, 8'd164, 8'd120, 8'd151, 8'd134, 8'd139, 8'd139, 8'd185, 8'd138, 8'd99, 8'd166, 8'd169, 8'd132, 8'd158, 8'd143, 8'd88, 8'd143, 8'd81, 8'd169, 8'd179, 8'd108, 8'd140, 8'd169, 8'd125, 8'd85, 8'd94, 8'd97, 8'd103, 8'd129, 8'd140, 8'd140, 8'd131, 8'd110, 8'd157, 8'd161, 8'd134, 8'd88, 8'd103, 8'd161, 8'd151, 8'd86, 8'd122, 8'd156, 8'd148, 8'd105, 8'd158, 8'd136, 8'd116, 8'd126, 8'd85, 8'd92, 8'd112, 8'd65, 8'd105, 8'd68, 8'd97, 8'd66, 8'd90, 8'd77, 8'd97, 8'd109, 8'd119, 8'd162, 8'd105, 8'd161, 8'd145, 8'd80, 8'd121, 8'd99, 8'd93, 8'd88, 8'd145, 8'd104, 8'd191, 8'd140, 8'd92, 8'd106, 8'd139, 8'd79, 8'd51, 8'd85, 8'd47, 8'd100, 8'd104, 8'd144, 8'd112, 8'd121, 8'd142, 8'd115, 8'd109, 8'd101, 8'd137, 8'd151, 8'd135, 8'd96, 8'd107, 8'd137, 8'd89, 8'd161, 8'd164, 8'd172, 8'd196, 8'd167, 8'd157, 8'd149, 8'd93, 8'd123, 8'd94, 8'd101, 8'd56, 8'd136, 8'd102, 8'd130, 8'd151, 8'd156, 8'd86, 8'd94, 8'd131, 8'd139, 8'd173, 8'd113, 8'd130, 8'd131, 8'd95, 8'd154, 8'd120, 8'd107, 8'd147, 8'd125, 8'd155, 8'd185, 8'd156, 8'd173, 8'd166, 8'd157, 8'd109, 8'd73, 8'd107, 8'd73, 8'd96, 8'd164, 8'd69, 8'd103, 8'd91, 8'd149, 8'd87, 8'd110, 8'd174, 8'd101, 8'd162, 8'd98, 8'd129, 8'd148, 8'd128, 8'd131, 8'd93, 8'd150, 8'd139, 8'd105, 8'd143, 8'd131, 8'd92, 8'd150, 8'd139, 8'd110, 8'd95, 8'd113, 8'd49, 8'd97, 8'd129, 8'd68, 8'd119, 8'd57, 8'd160, 8'd136, 8'd179, 8'd131, 8'd87, 8'd152, 8'd102, 8'd101, 8'd165, 8'd139, 8'd89, 8'd135, 8'd67, 8'd162, 8'd194, 8'd160, 8'd128, 8'd175, 8'd136, 8'd92, 8'd102, 8'd79, 8'd65, 8'd56, 8'd120, 8'd146, 8'd83, 8'd80, 8'd94, 8'd96, 8'd105, 8'd93, 8'd78, 8'd175, 8'd142, 8'd134, 8'd154, 8'd105, 8'd75, 8'd97, 8'd151, 8'd135, 8'd169, 8'd171, 8'd111, 8'd123, 8'd178, 8'd96, 8'd62, 8'd78, 8'd138, 8'd72, 8'd124, 8'd101, 8'd79, 8'd48, 8'd147, 8'd154, 8'd86, 8'd143, 8'd146, 8'd160, 8'd155, 8'd87, 8'd162, 8'd162, 8'd131, 8'd147, 8'd70, 8'd188, 8'd126, 8'd113, 8'd116, 8'd92, 8'd157, 8'd101, 8'd88, 8'd124, 8'd107, 8'd134, 8'd126, 8'd68, 8'd119, 8'd54, 8'd79, 8'd186, 8'd134, 8'd100, 8'd92, 8'd137, 8'd94, 8'd83, 8'd162, 8'd171, 8'd148, 8'd149, 8'd96, 8'd134, 8'd165, 8'd206, 8'd96, 8'd154, 8'd151, 8'd157, 8'd94, 8'd56, 8'd122, 8'd113, 8'd106, 8'd135, 8'd106, 8'd48, 8'd108, 8'd97, 8'd129, 8'd121, 8'd121, 8'd112, 8'd116, 8'd112, 8'd138, 8'd115, 8'd91, 8'd147, 8'd166, 8'd112, 8'd178, 8'd203, 8'd152, 8'd170, 8'd86, 8'd79, 8'd144, 8'd103, 8'd136, 8'd74, 8'd96, 8'd152, 8'd111, 8'd126, 8'd101, 8'd169, 8'd177, 8'd126, 8'd106, 8'd175, 8'd97, 8'd153, 8'd165, 8'd174, 8'd114, 8'd114, 8'd118, 8'd209, 8'd141, 8'd192, 8'd127, 8'd162, 8'd137, 8'd140, 8'd126, 8'd164, 8'd132, 8'd99, 8'd103, 8'd144, 8'd67, 8'd93, 8'd123, 8'd155, 8'd175, 8'd149, 8'd131, 8'd118, 8'd136, 8'd119, 8'd82, 8'd150, 8'd96, 8'd130, 8'd118, 8'd189, 8'd131, 8'd151, 8'd161, 8'd136, 8'd175, 8'd182, 8'd91, 8'd106, 8'd71, 8'd61, 8'd103, 8'd93, 8'd156, 8'd142, 8'd194, 8'd183, 8'd143, 8'd98, 8'd159, 8'd119, 8'd131, 8'd119, 8'd148, 8'd101, 8'd63, 8'd64, 8'd123, 8'd138, 8'd127, 8'd99, 8'd115, 8'd117, 8'd105, 8'd166, 8'd151, 8'd157, 8'd45, 8'd56, 8'd76, 8'd163, 8'd64, 8'd112, 8'd188, 8'd218, 8'd130, 8'd84, 8'd115, 8'd69, 8'd124, 8'd57, 8'd110, 8'd88, 8'd71, 8'd55, 8'd133, 8'd115, 8'd188, 8'd135, 8'd129, 8'd194, 8'd106, 8'd178, 8'd147, 8'd95, 8'd88, 8'd82, 8'd63, 8'd99, 8'd163, 8'd149, 8'd210, 8'd168, 8'd192, 8'd96, 8'd150, 8'd99, 8'd133, 8'd44, 8'd98, 8'd81, 8'd44, 8'd92, 8'd86, 8'd123, 8'd112, 8'd156, 8'd115, 8'd184, 8'd161, 8'd84, 8'd121, 8'd62, 8'd50, 8'd92, 8'd56, 8'd131, 8'd138, 8'd178, 8'd119, 8'd217, 8'd165, 8'd132, 8'd96, 8'd106, 8'd150, 8'd100, 8'd111, 8'd125, 8'd158, 8'd81, 8'd135, 8'd161, 8'd116, 8'd174, 8'd175, 8'd181, 8'd87, 8'd67, 8'd71, 8'd64, 8'd105, 8'd88, 8'd149, 8'd165, 8'd108, 8'd150, 8'd184, 8'd177, 8'd125, 8'd95, 8'd66, 8'd144, 8'd88, 8'd140, 8'd108, 8'd154, 8'd187, 8'd97, 8'd106, 8'd174, 8'd151, 8'd141, 8'd170, 8'd158, 8'd114, 8'd127, 8'd50, 8'd124, 8'd46, 8'd105, 8'd86, 8'd106, 8'd164, 8'd134, 8'd151, 8'd141, 8'd153, 8'd93, 8'd78, 8'd120, 8'd162, 8'd120, 8'd134, 8'd115, 8'd142, 8'd184, 8'd109, 8'd137, 8'd116, 8'd159, 8'd132, 8'd164, 8'd118, 8'd125, 8'd99, 8'd130, 8'd61, 8'd124, 8'd149, 8'd127, 8'd136, 8'd121, 8'd134, 8'd84, 8'd140, 8'd134, 8'd131, 8'd112, 8'd121, 8'd100, 8'd77, 8'd134, 8'd113, 8'd162, 8'd155, 8'd98, 8'd136, 8'd87, 8'd107, 8'd169, 8'd67, 8'd106, 8'd44, 8'd128, 8'd106, 8'd147, 8'd71, 8'd149, 8'd95, 8'd92, 8'd188, 8'd111, 8'd107, 8'd124, 8'd83, 8'd132, 8'd154, 8'd176, 8'd143, 8'd121, 8'd160, 8'd103, 8'd88, 8'd89, 8'd150, 8'd79, 8'd98, 8'd97, 8'd78, 8'd121, 8'd95, 8'd118, 8'd59, 8'd159, 8'd132, 8'd97, 8'd92, 8'd86, 8'd137, 8'd113, 8'd172, 8'd126, 8'd214, 8'd208, 8'd126, 8'd161, 8'd146, 8'd101, 8'd171, 8'd167, 8'd125, 8'd141, 8'd137, 8'd121, 8'd194, 8'd142, 8'd132, 8'd100, 8'd152, 8'd108, 8'd119, 8'd135, 8'd85, 8'd100, 8'd133, 8'd117, 8'd135, 8'd131, 8'd97, 8'd156, 8'd176, 8'd189, 8'd118, 8'd171, 8'd151, 8'd157, 8'd108, 8'd103, 8'd149, 8'd143, 8'd127, 8'd174, 8'd158, 8'd203, 8'd173, 8'd135, 8'd88, 8'd109, 8'd131, 8'd98, 8'd140, 8'd151, 8'd78, 8'd162, 8'd83, 8'd87, 8'd91, 8'd110, 8'd164, 8'd172, 8'd90, 8'd129, 8'd103, 8'd109, 8'd86, 8'd97, 8'd115, 8'd162, 8'd197, 8'd153, 8'd99, 8'd117, 8'd181, 8'd154, 8'd168, 8'd75, 8'd156, 8'd71, 8'd82, 8'd123, 8'd87, 8'd132, 8'd128, 8'd103, 8'd99, 8'd162, 8'd128, 8'd142, 8'd164, 8'd82, 8'd133, 8'd80, 8'd163, 8'd152, 8'd144, 8'd145, 8'd161, 8'd78, 8'd93, 8'd106, 8'd138, 8'd100, 8'd77, 8'd154, 8'd72, 8'd97, 8'd151, 8'd97})
) cell_0_66 (
    .clk(clk),
    .input_index(index_0_65_66),
    .input_value(value_0_65_66),
    .input_result(result_0_65_66),
    .input_enable(enable_0_65_66),
    .output_index(index_0_66_67),
    .output_value(value_0_66_67),
    .output_result(result_0_66_67),
    .output_enable(enable_0_66_67)
);

wire [10-1:0] index_0_67_68;
wire [`DATA_WIDTH-1:0] value_0_67_68;
wire [`DATA_WIDTH*4:0] result_0_67_68;
wire enable_0_67_68;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd142, 8'd97, 8'd102, 8'd165, 8'd126, 8'd84, 8'd159, 8'd105, 8'd157, 8'd127, 8'd205, 8'd194, 8'd100, 8'd132, 8'd157, 8'd125, 8'd78, 8'd134, 8'd106, 8'd137, 8'd142, 8'd162, 8'd101, 8'd168, 8'd164, 8'd106, 8'd93, 8'd114, 8'd162, 8'd123, 8'd109, 8'd109, 8'd83, 8'd170, 8'd120, 8'd124, 8'd131, 8'd140, 8'd114, 8'd105, 8'd112, 8'd148, 8'd119, 8'd127, 8'd99, 8'd107, 8'd89, 8'd175, 8'd111, 8'd99, 8'd110, 8'd129, 8'd147, 8'd70, 8'd73, 8'd93, 8'd160, 8'd97, 8'd128, 8'd80, 8'd137, 8'd75, 8'd96, 8'd161, 8'd107, 8'd147, 8'd125, 8'd170, 8'd118, 8'd97, 8'd148, 8'd148, 8'd149, 8'd126, 8'd97, 8'd165, 8'd149, 8'd121, 8'd182, 8'd174, 8'd108, 8'd153, 8'd85, 8'd87, 8'd130, 8'd94, 8'd150, 8'd143, 8'd74, 8'd77, 8'd150, 8'd64, 8'd84, 8'd78, 8'd123, 8'd93, 8'd118, 8'd110, 8'd143, 8'd144, 8'd91, 8'd103, 8'd113, 8'd72, 8'd76, 8'd114, 8'd116, 8'd150, 8'd110, 8'd83, 8'd127, 8'd75, 8'd80, 8'd68, 8'd131, 8'd146, 8'd131, 8'd161, 8'd89, 8'd122, 8'd89, 8'd130, 8'd76, 8'd113, 8'd82, 8'd113, 8'd139, 8'd100, 8'd122, 8'd108, 8'd114, 8'd69, 8'd133, 8'd105, 8'd67, 8'd46, 8'd44, 8'd126, 8'd128, 8'd161, 8'd137, 8'd153, 8'd71, 8'd145, 8'd87, 8'd154, 8'd67, 8'd133, 8'd121, 8'd100, 8'd96, 8'd91, 8'd136, 8'd152, 8'd173, 8'd131, 8'd168, 8'd154, 8'd84, 8'd100, 8'd107, 8'd152, 8'd84, 8'd81, 8'd116, 8'd97, 8'd155, 8'd109, 8'd160, 8'd125, 8'd160, 8'd165, 8'd121, 8'd60, 8'd130, 8'd48, 8'd100, 8'd109, 8'd146, 8'd121, 8'd101, 8'd148, 8'd113, 8'd149, 8'd167, 8'd140, 8'd106, 8'd82, 8'd128, 8'd118, 8'd92, 8'd86, 8'd67, 8'd136, 8'd81, 8'd68, 8'd66, 8'd169, 8'd107, 8'd109, 8'd65, 8'd119, 8'd116, 8'd87, 8'd78, 8'd61, 8'd137, 8'd131, 8'd119, 8'd138, 8'd120, 8'd186, 8'd134, 8'd79, 8'd106, 8'd145, 8'd140, 8'd112, 8'd121, 8'd87, 8'd52, 8'd152, 8'd168, 8'd73, 8'd148, 8'd122, 8'd126, 8'd92, 8'd87, 8'd115, 8'd122, 8'd83, 8'd94, 8'd100, 8'd144, 8'd128, 8'd160, 8'd121, 8'd168, 8'd188, 8'd189, 8'd112, 8'd158, 8'd125, 8'd126, 8'd107, 8'd78, 8'd119, 8'd31, 8'd157, 8'd166, 8'd87, 8'd109, 8'd73, 8'd147, 8'd166, 8'd148, 8'd106, 8'd130, 8'd92, 8'd91, 8'd144, 8'd99, 8'd167, 8'd111, 8'd156, 8'd95, 8'd160, 8'd123, 8'd108, 8'd165, 8'd117, 8'd111, 8'd160, 8'd134, 8'd108, 8'd90, 8'd128, 8'd155, 8'd162, 8'd108, 8'd97, 8'd96, 8'd99, 8'd98, 8'd70, 8'd164, 8'd78, 8'd83, 8'd161, 8'd85, 8'd168, 8'd102, 8'd107, 8'd123, 8'd104, 8'd144, 8'd122, 8'd117, 8'd136, 8'd137, 8'd97, 8'd158, 8'd111, 8'd107, 8'd140, 8'd92, 8'd121, 8'd91, 8'd71, 8'd143, 8'd77, 8'd110, 8'd148, 8'd125, 8'd108, 8'd164, 8'd99, 8'd89, 8'd111, 8'd115, 8'd72, 8'd60, 8'd81, 8'd108, 8'd129, 8'd158, 8'd184, 8'd155, 8'd188, 8'd129, 8'd155, 8'd59, 8'd84, 8'd125, 8'd158, 8'd149, 8'd131, 8'd108, 8'd160, 8'd138, 8'd121, 8'd177, 8'd155, 8'd89, 8'd153, 8'd167, 8'd156, 8'd88, 8'd67, 8'd94, 8'd77, 8'd80, 8'd188, 8'd168, 8'd177, 8'd156, 8'd165, 8'd154, 8'd127, 8'd146, 8'd72, 8'd88, 8'd151, 8'd92, 8'd95, 8'd131, 8'd183, 8'd125, 8'd162, 8'd163, 8'd154, 8'd142, 8'd161, 8'd92, 8'd108, 8'd114, 8'd46, 8'd97, 8'd135, 8'd161, 8'd110, 8'd125, 8'd119, 8'd107, 8'd178, 8'd136, 8'd133, 8'd75, 8'd115, 8'd107, 8'd67, 8'd80, 8'd71, 8'd132, 8'd184, 8'd165, 8'd174, 8'd168, 8'd172, 8'd155, 8'd159, 8'd142, 8'd95, 8'd34, 8'd29, 8'd66, 8'd119, 8'd120, 8'd114, 8'd174, 8'd139, 8'd147, 8'd164, 8'd148, 8'd132, 8'd108, 8'd132, 8'd124, 8'd142, 8'd164, 8'd68, 8'd103, 8'd127, 8'd143, 8'd145, 8'd123, 8'd105, 8'd114, 8'd111, 8'd166, 8'd106, 8'd28, 8'd31, 8'd39, 8'd96, 8'd150, 8'd153, 8'd165, 8'd89, 8'd103, 8'd111, 8'd137, 8'd77, 8'd113, 8'd128, 8'd145, 8'd149, 8'd122, 8'd70, 8'd88, 8'd109, 8'd172, 8'd103, 8'd120, 8'd151, 8'd134, 8'd128, 8'd167, 8'd96, 8'd40, 8'd130, 8'd109, 8'd149, 8'd169, 8'd108, 8'd154, 8'd137, 8'd165, 8'd140, 8'd111, 8'd98, 8'd164, 8'd116, 8'd177, 8'd92, 8'd113, 8'd118, 8'd32, 8'd114, 8'd140, 8'd137, 8'd145, 8'd145, 8'd104, 8'd128, 8'd157, 8'd119, 8'd83, 8'd116, 8'd101, 8'd150, 8'd167, 8'd163, 8'd144, 8'd138, 8'd157, 8'd91, 8'd83, 8'd110, 8'd160, 8'd148, 8'd103, 8'd123, 8'd73, 8'd101, 8'd88, 8'd53, 8'd124, 8'd120, 8'd120, 8'd116, 8'd166, 8'd126, 8'd183, 8'd107, 8'd97, 8'd119, 8'd119, 8'd118, 8'd157, 8'd82, 8'd164, 8'd125, 8'd94, 8'd115, 8'd155, 8'd83, 8'd98, 8'd96, 8'd89, 8'd158, 8'd146, 8'd64, 8'd71, 8'd106, 8'd132, 8'd153, 8'd103, 8'd121, 8'd142, 8'd174, 8'd151, 8'd149, 8'd112, 8'd109, 8'd122, 8'd156, 8'd137, 8'd158, 8'd178, 8'd98, 8'd86, 8'd111, 8'd168, 8'd105, 8'd142, 8'd168, 8'd97, 8'd115, 8'd106, 8'd86, 8'd86, 8'd102, 8'd131, 8'd137, 8'd89, 8'd90, 8'd160, 8'd129, 8'd161, 8'd144, 8'd142, 8'd87, 8'd91, 8'd79, 8'd96, 8'd123, 8'd101, 8'd120, 8'd104, 8'd80, 8'd105, 8'd113, 8'd157, 8'd129, 8'd154, 8'd135, 8'd158, 8'd97, 8'd97, 8'd75, 8'd99, 8'd96, 8'd105, 8'd83, 8'd109, 8'd133, 8'd118, 8'd138, 8'd147, 8'd80, 8'd138, 8'd102, 8'd89, 8'd79, 8'd78, 8'd171, 8'd80, 8'd150, 8'd122, 8'd143, 8'd82, 8'd161, 8'd147, 8'd149, 8'd157, 8'd84, 8'd56, 8'd68, 8'd134, 8'd160, 8'd140, 8'd137, 8'd69, 8'd123, 8'd82, 8'd150, 8'd159, 8'd65, 8'd99, 8'd132, 8'd150, 8'd105, 8'd101, 8'd169, 8'd83, 8'd118, 8'd119, 8'd116, 8'd101, 8'd69, 8'd131, 8'd80, 8'd152, 8'd163, 8'd139, 8'd75, 8'd98, 8'd172, 8'd72, 8'd105, 8'd107, 8'd122, 8'd162, 8'd118, 8'd136, 8'd116, 8'd126, 8'd90, 8'd59, 8'd94, 8'd113, 8'd139, 8'd149, 8'd117, 8'd140, 8'd118, 8'd98, 8'd84, 8'd156, 8'd138, 8'd141, 8'd102, 8'd149, 8'd174, 8'd114, 8'd175, 8'd170, 8'd73, 8'd94, 8'd96, 8'd90, 8'd139, 8'd116, 8'd156, 8'd131, 8'd159, 8'd101, 8'd108, 8'd165, 8'd105, 8'd117, 8'd86, 8'd94, 8'd157, 8'd90, 8'd87, 8'd74, 8'd140, 8'd104, 8'd125, 8'd129, 8'd82, 8'd135, 8'd126, 8'd149, 8'd133, 8'd153, 8'd96, 8'd112, 8'd130, 8'd124, 8'd180, 8'd135, 8'd130, 8'd141, 8'd195, 8'd121, 8'd127, 8'd147, 8'd131, 8'd109, 8'd81, 8'd83, 8'd126, 8'd162, 8'd161, 8'd157, 8'd143, 8'd93, 8'd96, 8'd139, 8'd159, 8'd117, 8'd163, 8'd150, 8'd133, 8'd165, 8'd181, 8'd125, 8'd168, 8'd126, 8'd175, 8'd153, 8'd177, 8'd148, 8'd109, 8'd117, 8'd96, 8'd121, 8'd150, 8'd161, 8'd111, 8'd117, 8'd94, 8'd114, 8'd80, 8'd132, 8'd109, 8'd117, 8'd142, 8'd79, 8'd80, 8'd114, 8'd137, 8'd99, 8'd125, 8'd132, 8'd71, 8'd147, 8'd113, 8'd113, 8'd105, 8'd87, 8'd80, 8'd129, 8'd97, 8'd167, 8'd150, 8'd147, 8'd163, 8'd89, 8'd129})
) cell_0_67 (
    .clk(clk),
    .input_index(index_0_66_67),
    .input_value(value_0_66_67),
    .input_result(result_0_66_67),
    .input_enable(enable_0_66_67),
    .output_index(index_0_67_68),
    .output_value(value_0_67_68),
    .output_result(result_0_67_68),
    .output_enable(enable_0_67_68)
);

wire [10-1:0] index_0_68_69;
wire [`DATA_WIDTH-1:0] value_0_68_69;
wire [`DATA_WIDTH*4:0] result_0_68_69;
wire enable_0_68_69;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd170, 8'd104, 8'd79, 8'd114, 8'd110, 8'd173, 8'd135, 8'd170, 8'd137, 8'd128, 8'd175, 8'd88, 8'd114, 8'd111, 8'd152, 8'd141, 8'd123, 8'd67, 8'd89, 8'd95, 8'd143, 8'd151, 8'd104, 8'd148, 8'd138, 8'd85, 8'd79, 8'd114, 8'd79, 8'd119, 8'd87, 8'd92, 8'd69, 8'd97, 8'd83, 8'd49, 8'd95, 8'd86, 8'd117, 8'd33, 8'd111, 8'd68, 8'd76, 8'd114, 8'd63, 8'd103, 8'd115, 8'd80, 8'd62, 8'd90, 8'd149, 8'd87, 8'd101, 8'd88, 8'd166, 8'd166, 8'd70, 8'd176, 8'd153, 8'd142, 8'd145, 8'd123, 8'd115, 8'd53, 8'd42, 8'd74, 8'd115, 8'd102, 8'd103, 8'd128, 8'd77, 8'd69, 8'd44, 8'd121, 8'd45, 8'd57, 8'd118, 8'd90, 8'd149, 8'd106, 8'd110, 8'd150, 8'd81, 8'd148, 8'd167, 8'd82, 8'd150, 8'd91, 8'd53, 8'd135, 8'd140, 8'd97, 8'd155, 8'd161, 8'd160, 8'd121, 8'd92, 8'd82, 8'd80, 8'd89, 8'd96, 8'd143, 8'd136, 8'd75, 8'd129, 8'd91, 8'd87, 8'd101, 8'd142, 8'd176, 8'd119, 8'd169, 8'd102, 8'd137, 8'd142, 8'd129, 8'd115, 8'd70, 8'd117, 8'd116, 8'd144, 8'd153, 8'd93, 8'd147, 8'd90, 8'd128, 8'd120, 8'd104, 8'd54, 8'd53, 8'd99, 8'd109, 8'd137, 8'd168, 8'd155, 8'd94, 8'd153, 8'd160, 8'd131, 8'd133, 8'd106, 8'd116, 8'd71, 8'd93, 8'd120, 8'd147, 8'd97, 8'd132, 8'd107, 8'd102, 8'd115, 8'd82, 8'd150, 8'd141, 8'd91, 8'd149, 8'd67, 8'd147, 8'd132, 8'd62, 8'd101, 8'd118, 8'd139, 8'd146, 8'd95, 8'd109, 8'd142, 8'd117, 8'd83, 8'd160, 8'd99, 8'd119, 8'd144, 8'd103, 8'd121, 8'd79, 8'd81, 8'd93, 8'd165, 8'd117, 8'd149, 8'd122, 8'd148, 8'd128, 8'd71, 8'd77, 8'd116, 8'd101, 8'd90, 8'd151, 8'd101, 8'd126, 8'd115, 8'd136, 8'd168, 8'd126, 8'd136, 8'd136, 8'd159, 8'd131, 8'd70, 8'd149, 8'd78, 8'd89, 8'd130, 8'd157, 8'd125, 8'd154, 8'd153, 8'd143, 8'd149, 8'd77, 8'd80, 8'd67, 8'd80, 8'd118, 8'd91, 8'd142, 8'd85, 8'd134, 8'd174, 8'd122, 8'd95, 8'd109, 8'd117, 8'd113, 8'd97, 8'd121, 8'd91, 8'd78, 8'd151, 8'd124, 8'd99, 8'd93, 8'd125, 8'd122, 8'd87, 8'd86, 8'd116, 8'd118, 8'd139, 8'd78, 8'd55, 8'd85, 8'd149, 8'd87, 8'd45, 8'd97, 8'd117, 8'd125, 8'd138, 8'd135, 8'd123, 8'd124, 8'd150, 8'd95, 8'd122, 8'd84, 8'd167, 8'd141, 8'd83, 8'd88, 8'd69, 8'd77, 8'd137, 8'd127, 8'd159, 8'd92, 8'd121, 8'd150, 8'd143, 8'd72, 8'd106, 8'd53, 8'd142, 8'd145, 8'd142, 8'd182, 8'd90, 8'd103, 8'd124, 8'd114, 8'd154, 8'd55, 8'd87, 8'd154, 8'd148, 8'd92, 8'd139, 8'd72, 8'd117, 8'd97, 8'd102, 8'd142, 8'd147, 8'd186, 8'd130, 8'd125, 8'd106, 8'd139, 8'd123, 8'd110, 8'd119, 8'd83, 8'd108, 8'd170, 8'd179, 8'd143, 8'd152, 8'd141, 8'd148, 8'd134, 8'd66, 8'd108, 8'd92, 8'd135, 8'd74, 8'd138, 8'd151, 8'd134, 8'd190, 8'd169, 8'd124, 8'd108, 8'd120, 8'd143, 8'd102, 8'd162, 8'd88, 8'd141, 8'd155, 8'd115, 8'd130, 8'd162, 8'd82, 8'd173, 8'd95, 8'd92, 8'd112, 8'd73, 8'd71, 8'd131, 8'd88, 8'd134, 8'd124, 8'd141, 8'd109, 8'd135, 8'd203, 8'd133, 8'd185, 8'd96, 8'd165, 8'd88, 8'd81, 8'd108, 8'd150, 8'd145, 8'd127, 8'd97, 8'd95, 8'd92, 8'd157, 8'd149, 8'd134, 8'd71, 8'd175, 8'd118, 8'd126, 8'd143, 8'd169, 8'd161, 8'd141, 8'd123, 8'd117, 8'd114, 8'd176, 8'd158, 8'd166, 8'd177, 8'd171, 8'd130, 8'd79, 8'd157, 8'd83, 8'd140, 8'd144, 8'd93, 8'd145, 8'd165, 8'd106, 8'd80, 8'd106, 8'd108, 8'd109, 8'd99, 8'd179, 8'd176, 8'd144, 8'd164, 8'd130, 8'd148, 8'd134, 8'd147, 8'd201, 8'd205, 8'd175, 8'd76, 8'd75, 8'd106, 8'd143, 8'd121, 8'd113, 8'd164, 8'd81, 8'd105, 8'd110, 8'd112, 8'd140, 8'd175, 8'd79, 8'd66, 8'd138, 8'd190, 8'd171, 8'd183, 8'd134, 8'd128, 8'd72, 8'd154, 8'd81, 8'd104, 8'd105, 8'd148, 8'd122, 8'd165, 8'd151, 8'd83, 8'd123, 8'd141, 8'd119, 8'd76, 8'd60, 8'd62, 8'd81, 8'd148, 8'd69, 8'd123, 8'd124, 8'd103, 8'd115, 8'd83, 8'd157, 8'd92, 8'd118, 8'd84, 8'd155, 8'd123, 8'd156, 8'd99, 8'd164, 8'd176, 8'd101, 8'd149, 8'd72, 8'd115, 8'd149, 8'd130, 8'd80, 8'd148, 8'd138, 8'd111, 8'd90, 8'd116, 8'd78, 8'd90, 8'd81, 8'd46, 8'd82, 8'd44, 8'd123, 8'd135, 8'd89, 8'd115, 8'd159, 8'd95, 8'd155, 8'd148, 8'd92, 8'd113, 8'd144, 8'd125, 8'd60, 8'd80, 8'd71, 8'd102, 8'd121, 8'd69, 8'd153, 8'd114, 8'd129, 8'd121, 8'd175, 8'd166, 8'd125, 8'd99, 8'd95, 8'd83, 8'd78, 8'd120, 8'd86, 8'd67, 8'd126, 8'd74, 8'd137, 8'd102, 8'd148, 8'd119, 8'd110, 8'd128, 8'd103, 8'd123, 8'd152, 8'd124, 8'd86, 8'd150, 8'd100, 8'd99, 8'd127, 8'd146, 8'd73, 8'd95, 8'd141, 8'd71, 8'd63, 8'd80, 8'd87, 8'd120, 8'd118, 8'd88, 8'd129, 8'd144, 8'd61, 8'd112, 8'd42, 8'd61, 8'd112, 8'd69, 8'd139, 8'd57, 8'd123, 8'd130, 8'd119, 8'd132, 8'd149, 8'd201, 8'd165, 8'd121, 8'd96, 8'd131, 8'd165, 8'd146, 8'd87, 8'd71, 8'd101, 8'd72, 8'd98, 8'd118, 8'd140, 8'd102, 8'd60, 8'd36, 8'd114, 8'd67, 8'd65, 8'd56, 8'd49, 8'd141, 8'd87, 8'd137, 8'd78, 8'd166, 8'd166, 8'd175, 8'd90, 8'd134, 8'd107, 8'd84, 8'd107, 8'd131, 8'd100, 8'd82, 8'd144, 8'd157, 8'd93, 8'd145, 8'd88, 8'd133, 8'd84, 8'd83, 8'd82, 8'd118, 8'd150, 8'd63, 8'd67, 8'd120, 8'd146, 8'd134, 8'd124, 8'd176, 8'd156, 8'd188, 8'd127, 8'd118, 8'd153, 8'd105, 8'd171, 8'd88, 8'd99, 8'd135, 8'd133, 8'd132, 8'd138, 8'd95, 8'd118, 8'd130, 8'd105, 8'd96, 8'd108, 8'd96, 8'd81, 8'd71, 8'd121, 8'd93, 8'd101, 8'd165, 8'd99, 8'd143, 8'd123, 8'd160, 8'd134, 8'd88, 8'd99, 8'd83, 8'd85, 8'd94, 8'd91, 8'd76, 8'd162, 8'd170, 8'd102, 8'd193, 8'd148, 8'd77, 8'd111, 8'd99, 8'd160, 8'd96, 8'd92, 8'd133, 8'd127, 8'd82, 8'd111, 8'd98, 8'd178, 8'd172, 8'd136, 8'd164, 8'd97, 8'd157, 8'd171, 8'd80, 8'd102, 8'd99, 8'd171, 8'd159, 8'd94, 8'd148, 8'd94, 8'd94, 8'd152, 8'd83, 8'd140, 8'd118, 8'd140, 8'd137, 8'd143, 8'd127, 8'd88, 8'd89, 8'd100, 8'd136, 8'd157, 8'd133, 8'd110, 8'd126, 8'd81, 8'd134, 8'd87, 8'd80, 8'd112, 8'd83, 8'd137, 8'd160, 8'd144, 8'd114, 8'd163, 8'd135, 8'd88, 8'd97, 8'd142, 8'd129, 8'd168, 8'd167, 8'd124, 8'd105, 8'd117, 8'd164, 8'd99, 8'd115, 8'd138, 8'd87, 8'd131, 8'd85, 8'd155, 8'd169, 8'd81, 8'd97, 8'd81, 8'd105, 8'd135, 8'd81, 8'd124, 8'd78, 8'd155, 8'd116, 8'd109, 8'd103, 8'd98, 8'd66, 8'd90, 8'd95, 8'd119, 8'd155, 8'd145, 8'd62, 8'd110, 8'd109, 8'd94, 8'd62, 8'd155, 8'd155, 8'd127, 8'd151, 8'd104, 8'd92, 8'd132, 8'd108, 8'd84, 8'd105, 8'd125, 8'd72, 8'd149, 8'd137, 8'd160, 8'd100, 8'd88, 8'd131, 8'd82, 8'd164, 8'd117, 8'd129, 8'd99, 8'd81, 8'd157, 8'd156, 8'd105, 8'd122, 8'd116, 8'd142, 8'd134, 8'd152, 8'd104, 8'd165})
) cell_0_68 (
    .clk(clk),
    .input_index(index_0_67_68),
    .input_value(value_0_67_68),
    .input_result(result_0_67_68),
    .input_enable(enable_0_67_68),
    .output_index(index_0_68_69),
    .output_value(value_0_68_69),
    .output_result(result_0_68_69),
    .output_enable(enable_0_68_69)
);

wire [10-1:0] index_0_69_70;
wire [`DATA_WIDTH-1:0] value_0_69_70;
wire [`DATA_WIDTH*4:0] result_0_69_70;
wire enable_0_69_70;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd167, 8'd113, 8'd120, 8'd154, 8'd178, 8'd72, 8'd160, 8'd145, 8'd83, 8'd93, 8'd88, 8'd100, 8'd103, 8'd150, 8'd138, 8'd162, 8'd131, 8'd167, 8'd137, 8'd91, 8'd135, 8'd134, 8'd77, 8'd133, 8'd160, 8'd97, 8'd125, 8'd151, 8'd169, 8'd117, 8'd155, 8'd108, 8'd123, 8'd130, 8'd144, 8'd96, 8'd63, 8'd138, 8'd130, 8'd61, 8'd146, 8'd111, 8'd111, 8'd70, 8'd77, 8'd141, 8'd133, 8'd51, 8'd120, 8'd127, 8'd125, 8'd98, 8'd127, 8'd116, 8'd72, 8'd125, 8'd167, 8'd155, 8'd165, 8'd109, 8'd167, 8'd140, 8'd122, 8'd144, 8'd98, 8'd154, 8'd131, 8'd123, 8'd155, 8'd98, 8'd140, 8'd118, 8'd141, 8'd102, 8'd132, 8'd53, 8'd67, 8'd78, 8'd102, 8'd75, 8'd137, 8'd157, 8'd88, 8'd81, 8'd136, 8'd155, 8'd88, 8'd176, 8'd113, 8'd125, 8'd157, 8'd163, 8'd98, 8'd146, 8'd124, 8'd169, 8'd145, 8'd109, 8'd121, 8'd135, 8'd146, 8'd136, 8'd116, 8'd132, 8'd71, 8'd76, 8'd81, 8'd125, 8'd90, 8'd86, 8'd97, 8'd146, 8'd94, 8'd155, 8'd158, 8'd176, 8'd98, 8'd149, 8'd111, 8'd130, 8'd162, 8'd114, 8'd146, 8'd152, 8'd147, 8'd103, 8'd177, 8'd158, 8'd122, 8'd128, 8'd133, 8'd141, 8'd122, 8'd74, 8'd67, 8'd163, 8'd138, 8'd102, 8'd98, 8'd79, 8'd165, 8'd101, 8'd111, 8'd120, 8'd102, 8'd179, 8'd101, 8'd110, 8'd170, 8'd101, 8'd109, 8'd140, 8'd127, 8'd135, 8'd88, 8'd153, 8'd116, 8'd74, 8'd101, 8'd142, 8'd94, 8'd106, 8'd100, 8'd90, 8'd93, 8'd107, 8'd75, 8'd78, 8'd81, 8'd115, 8'd162, 8'd175, 8'd186, 8'd190, 8'd94, 8'd117, 8'd66, 8'd150, 8'd77, 8'd121, 8'd88, 8'd132, 8'd111, 8'd81, 8'd74, 8'd110, 8'd147, 8'd103, 8'd152, 8'd143, 8'd144, 8'd129, 8'd94, 8'd149, 8'd141, 8'd93, 8'd128, 8'd116, 8'd156, 8'd131, 8'd182, 8'd149, 8'd117, 8'd114, 8'd69, 8'd123, 8'd69, 8'd68, 8'd152, 8'd102, 8'd90, 8'd127, 8'd75, 8'd138, 8'd77, 8'd121, 8'd92, 8'd138, 8'd102, 8'd157, 8'd56, 8'd163, 8'd123, 8'd103, 8'd75, 8'd132, 8'd92, 8'd160, 8'd137, 8'd132, 8'd153, 8'd94, 8'd95, 8'd111, 8'd113, 8'd81, 8'd148, 8'd144, 8'd137, 8'd150, 8'd150, 8'd75, 8'd83, 8'd81, 8'd159, 8'd156, 8'd160, 8'd116, 8'd74, 8'd93, 8'd73, 8'd113, 8'd88, 8'd172, 8'd65, 8'd114, 8'd110, 8'd97, 8'd148, 8'd102, 8'd95, 8'd84, 8'd78, 8'd157, 8'd158, 8'd127, 8'd108, 8'd107, 8'd102, 8'd121, 8'd148, 8'd117, 8'd111, 8'd139, 8'd88, 8'd150, 8'd107, 8'd70, 8'd93, 8'd157, 8'd148, 8'd166, 8'd131, 8'd120, 8'd133, 8'd98, 8'd135, 8'd118, 8'd95, 8'd140, 8'd80, 8'd118, 8'd166, 8'd178, 8'd145, 8'd95, 8'd82, 8'd162, 8'd117, 8'd130, 8'd157, 8'd117, 8'd154, 8'd105, 8'd49, 8'd134, 8'd63, 8'd166, 8'd129, 8'd164, 8'd62, 8'd106, 8'd156, 8'd63, 8'd90, 8'd66, 8'd86, 8'd89, 8'd166, 8'd178, 8'd167, 8'd71, 8'd85, 8'd87, 8'd167, 8'd113, 8'd82, 8'd80, 8'd159, 8'd81, 8'd120, 8'd79, 8'd84, 8'd73, 8'd92, 8'd135, 8'd123, 8'd166, 8'd130, 8'd112, 8'd124, 8'd107, 8'd122, 8'd126, 8'd112, 8'd92, 8'd94, 8'd160, 8'd83, 8'd101, 8'd140, 8'd91, 8'd80, 8'd141, 8'd78, 8'd168, 8'd137, 8'd118, 8'd101, 8'd174, 8'd157, 8'd112, 8'd113, 8'd161, 8'd78, 8'd144, 8'd73, 8'd132, 8'd76, 8'd163, 8'd117, 8'd77, 8'd85, 8'd99, 8'd149, 8'd133, 8'd83, 8'd130, 8'd138, 8'd167, 8'd142, 8'd100, 8'd137, 8'd110, 8'd97, 8'd173, 8'd133, 8'd159, 8'd157, 8'd70, 8'd91, 8'd145, 8'd139, 8'd139, 8'd75, 8'd130, 8'd91, 8'd102, 8'd111, 8'd95, 8'd89, 8'd78, 8'd54, 8'd63, 8'd71, 8'd106, 8'd62, 8'd151, 8'd107, 8'd170, 8'd164, 8'd142, 8'd157, 8'd183, 8'd174, 8'd98, 8'd138, 8'd143, 8'd164, 8'd96, 8'd146, 8'd158, 8'd87, 8'd79, 8'd102, 8'd72, 8'd140, 8'd73, 8'd67, 8'd119, 8'd123, 8'd148, 8'd80, 8'd100, 8'd91, 8'd155, 8'd177, 8'd88, 8'd171, 8'd168, 8'd126, 8'd143, 8'd169, 8'd139, 8'd69, 8'd80, 8'd75, 8'd88, 8'd146, 8'd161, 8'd162, 8'd100, 8'd89, 8'd92, 8'd131, 8'd95, 8'd147, 8'd68, 8'd130, 8'd124, 8'd90, 8'd67, 8'd134, 8'd125, 8'd156, 8'd148, 8'd191, 8'd201, 8'd165, 8'd179, 8'd163, 8'd105, 8'd114, 8'd57, 8'd145, 8'd100, 8'd104, 8'd182, 8'd143, 8'd226, 8'd145, 8'd134, 8'd181, 8'd139, 8'd154, 8'd105, 8'd124, 8'd134, 8'd130, 8'd91, 8'd142, 8'd161, 8'd161, 8'd189, 8'd180, 8'd156, 8'd180, 8'd98, 8'd162, 8'd122, 8'd62, 8'd140, 8'd90, 8'd137, 8'd86, 8'd140, 8'd220, 8'd194, 8'd127, 8'd197, 8'd140, 8'd130, 8'd137, 8'd153, 8'd90, 8'd113, 8'd129, 8'd75, 8'd73, 8'd139, 8'd181, 8'd150, 8'd145, 8'd117, 8'd150, 8'd161, 8'd120, 8'd75, 8'd70, 8'd108, 8'd120, 8'd80, 8'd147, 8'd120, 8'd180, 8'd204, 8'd212, 8'd180, 8'd152, 8'd102, 8'd101, 8'd133, 8'd127, 8'd90, 8'd127, 8'd101, 8'd115, 8'd144, 8'd157, 8'd79, 8'd154, 8'd152, 8'd135, 8'd74, 8'd125, 8'd103, 8'd66, 8'd172, 8'd94, 8'd139, 8'd143, 8'd134, 8'd148, 8'd207, 8'd130, 8'd117, 8'd93, 8'd169, 8'd127, 8'd97, 8'd128, 8'd62, 8'd55, 8'd130, 8'd88, 8'd107, 8'd85, 8'd105, 8'd144, 8'd115, 8'd115, 8'd128, 8'd106, 8'd122, 8'd130, 8'd175, 8'd135, 8'd94, 8'd125, 8'd157, 8'd162, 8'd173, 8'd128, 8'd138, 8'd162, 8'd114, 8'd107, 8'd151, 8'd91, 8'd156, 8'd91, 8'd58, 8'd55, 8'd147, 8'd106, 8'd107, 8'd63, 8'd154, 8'd112, 8'd69, 8'd94, 8'd111, 8'd89, 8'd146, 8'd72, 8'd120, 8'd129, 8'd166, 8'd174, 8'd158, 8'd176, 8'd129, 8'd144, 8'd107, 8'd113, 8'd104, 8'd107, 8'd99, 8'd131, 8'd102, 8'd65, 8'd121, 8'd139, 8'd128, 8'd153, 8'd78, 8'd103, 8'd89, 8'd123, 8'd93, 8'd150, 8'd123, 8'd139, 8'd115, 8'd113, 8'd156, 8'd136, 8'd105, 8'd86, 8'd91, 8'd76, 8'd158, 8'd134, 8'd74, 8'd164, 8'd138, 8'd159, 8'd109, 8'd105, 8'd145, 8'd109, 8'd127, 8'd85, 8'd126, 8'd75, 8'd48, 8'd57, 8'd110, 8'd81, 8'd139, 8'd75, 8'd129, 8'd169, 8'd149, 8'd143, 8'd126, 8'd147, 8'd131, 8'd133, 8'd115, 8'd134, 8'd58, 8'd81, 8'd84, 8'd105, 8'd91, 8'd75, 8'd121, 8'd108, 8'd49, 8'd63, 8'd120, 8'd47, 8'd122, 8'd113, 8'd116, 8'd109, 8'd66, 8'd102, 8'd166, 8'd129, 8'd95, 8'd100, 8'd124, 8'd141, 8'd126, 8'd68, 8'd58, 8'd47, 8'd58, 8'd57, 8'd88, 8'd70, 8'd49, 8'd31, 8'd50, 8'd112, 8'd49, 8'd112, 8'd63, 8'd45, 8'd130, 8'd118, 8'd67, 8'd138, 8'd114, 8'd90, 8'd142, 8'd133, 8'd127, 8'd155, 8'd133, 8'd140, 8'd110, 8'd82, 8'd118, 8'd64, 8'd64, 8'd73, 8'd55, 8'd95, 8'd93, 8'd79, 8'd57, 8'd84, 8'd103, 8'd52, 8'd90, 8'd114, 8'd142, 8'd96, 8'd148, 8'd117, 8'd91, 8'd139, 8'd114, 8'd130, 8'd111, 8'd132, 8'd116, 8'd141, 8'd102, 8'd125, 8'd74, 8'd150, 8'd144, 8'd85, 8'd167, 8'd169, 8'd162, 8'd98, 8'd142, 8'd129, 8'd115, 8'd93, 8'd84, 8'd82, 8'd85, 8'd170, 8'd131, 8'd85, 8'd97, 8'd148, 8'd97})
) cell_0_69 (
    .clk(clk),
    .input_index(index_0_68_69),
    .input_value(value_0_68_69),
    .input_result(result_0_68_69),
    .input_enable(enable_0_68_69),
    .output_index(index_0_69_70),
    .output_value(value_0_69_70),
    .output_result(result_0_69_70),
    .output_enable(enable_0_69_70)
);

wire [10-1:0] index_0_70_71;
wire [`DATA_WIDTH-1:0] value_0_70_71;
wire [`DATA_WIDTH*4:0] result_0_70_71;
wire enable_0_70_71;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd169, 8'd129, 8'd131, 8'd129, 8'd128, 8'd61, 8'd68, 8'd94, 8'd132, 8'd138, 8'd80, 8'd49, 8'd137, 8'd43, 8'd63, 8'd154, 8'd154, 8'd135, 8'd127, 8'd98, 8'd62, 8'd62, 8'd87, 8'd77, 8'd95, 8'd154, 8'd119, 8'd99, 8'd151, 8'd89, 8'd69, 8'd74, 8'd66, 8'd81, 8'd133, 8'd154, 8'd49, 8'd66, 8'd49, 8'd58, 8'd73, 8'd45, 8'd96, 8'd125, 8'd57, 8'd87, 8'd77, 8'd94, 8'd98, 8'd89, 8'd146, 8'd88, 8'd169, 8'd160, 8'd85, 8'd146, 8'd148, 8'd98, 8'd130, 8'd134, 8'd99, 8'd64, 8'd69, 8'd142, 8'd128, 8'd151, 8'd73, 8'd129, 8'd98, 8'd93, 8'd171, 8'd79, 8'd178, 8'd117, 8'd83, 8'd151, 8'd112, 8'd91, 8'd78, 8'd98, 8'd81, 8'd115, 8'd118, 8'd70, 8'd126, 8'd95, 8'd156, 8'd98, 8'd98, 8'd100, 8'd101, 8'd175, 8'd112, 8'd188, 8'd97, 8'd150, 8'd138, 8'd152, 8'd153, 8'd178, 8'd119, 8'd108, 8'd145, 8'd99, 8'd170, 8'd129, 8'd82, 8'd99, 8'd90, 8'd92, 8'd160, 8'd117, 8'd92, 8'd120, 8'd84, 8'd125, 8'd133, 8'd100, 8'd135, 8'd107, 8'd123, 8'd199, 8'd169, 8'd92, 8'd124, 8'd156, 8'd177, 8'd185, 8'd157, 8'd150, 8'd166, 8'd142, 8'd137, 8'd164, 8'd101, 8'd139, 8'd151, 8'd136, 8'd95, 8'd108, 8'd125, 8'd105, 8'd127, 8'd102, 8'd111, 8'd190, 8'd122, 8'd143, 8'd176, 8'd99, 8'd167, 8'd83, 8'd74, 8'd94, 8'd149, 8'd103, 8'd115, 8'd91, 8'd102, 8'd147, 8'd127, 8'd168, 8'd113, 8'd148, 8'd148, 8'd145, 8'd96, 8'd106, 8'd85, 8'd114, 8'd93, 8'd86, 8'd97, 8'd95, 8'd171, 8'd143, 8'd162, 8'd115, 8'd143, 8'd157, 8'd96, 8'd139, 8'd89, 8'd81, 8'd82, 8'd155, 8'd138, 8'd153, 8'd168, 8'd153, 8'd170, 8'd145, 8'd167, 8'd161, 8'd147, 8'd153, 8'd109, 8'd90, 8'd156, 8'd171, 8'd151, 8'd106, 8'd171, 8'd132, 8'd171, 8'd155, 8'd89, 8'd167, 8'd155, 8'd117, 8'd66, 8'd75, 8'd64, 8'd117, 8'd145, 8'd132, 8'd172, 8'd140, 8'd154, 8'd193, 8'd202, 8'd180, 8'd141, 8'd112, 8'd117, 8'd115, 8'd134, 8'd97, 8'd155, 8'd160, 8'd122, 8'd109, 8'd151, 8'd110, 8'd98, 8'd92, 8'd125, 8'd67, 8'd102, 8'd106, 8'd115, 8'd106, 8'd81, 8'd146, 8'd196, 8'd197, 8'd207, 8'd170, 8'd122, 8'd162, 8'd64, 8'd146, 8'd111, 8'd145, 8'd169, 8'd170, 8'd141, 8'd177, 8'd135, 8'd108, 8'd101, 8'd89, 8'd114, 8'd126, 8'd174, 8'd146, 8'd94, 8'd118, 8'd46, 8'd61, 8'd143, 8'd78, 8'd115, 8'd147, 8'd105, 8'd205, 8'd182, 8'd149, 8'd131, 8'd97, 8'd99, 8'd121, 8'd166, 8'd95, 8'd160, 8'd165, 8'd152, 8'd82, 8'd150, 8'd109, 8'd103, 8'd188, 8'd91, 8'd71, 8'd72, 8'd157, 8'd113, 8'd142, 8'd122, 8'd80, 8'd84, 8'd84, 8'd140, 8'd138, 8'd136, 8'd159, 8'd83, 8'd104, 8'd165, 8'd211, 8'd176, 8'd101, 8'd108, 8'd135, 8'd121, 8'd75, 8'd149, 8'd115, 8'd190, 8'd93, 8'd149, 8'd73, 8'd128, 8'd156, 8'd154, 8'd79, 8'd116, 8'd63, 8'd109, 8'd91, 8'd144, 8'd122, 8'd102, 8'd155, 8'd161, 8'd155, 8'd134, 8'd134, 8'd113, 8'd158, 8'd102, 8'd84, 8'd76, 8'd89, 8'd171, 8'd108, 8'd103, 8'd92, 8'd121, 8'd162, 8'd164, 8'd165, 8'd145, 8'd94, 8'd101, 8'd111, 8'd135, 8'd75, 8'd133, 8'd178, 8'd143, 8'd145, 8'd125, 8'd112, 8'd134, 8'd114, 8'd115, 8'd69, 8'd81, 8'd84, 8'd95, 8'd80, 8'd87, 8'd131, 8'd151, 8'd102, 8'd117, 8'd174, 8'd146, 8'd190, 8'd138, 8'd155, 8'd153, 8'd86, 8'd117, 8'd145, 8'd60, 8'd74, 8'd97, 8'd127, 8'd159, 8'd132, 8'd147, 8'd147, 8'd133, 8'd67, 8'd121, 8'd114, 8'd67, 8'd117, 8'd165, 8'd121, 8'd184, 8'd100, 8'd85, 8'd180, 8'd182, 8'd142, 8'd146, 8'd124, 8'd125, 8'd59, 8'd41, 8'd70, 8'd92, 8'd72, 8'd142, 8'd63, 8'd64, 8'd108, 8'd122, 8'd136, 8'd138, 8'd74, 8'd82, 8'd58, 8'd93, 8'd133, 8'd152, 8'd103, 8'd140, 8'd97, 8'd100, 8'd172, 8'd84, 8'd136, 8'd108, 8'd166, 8'd104, 8'd130, 8'd113, 8'd81, 8'd76, 8'd111, 8'd123, 8'd72, 8'd125, 8'd141, 8'd120, 8'd158, 8'd175, 8'd91, 8'd97, 8'd137, 8'd134, 8'd150, 8'd134, 8'd124, 8'd102, 8'd101, 8'd122, 8'd123, 8'd114, 8'd71, 8'd98, 8'd56, 8'd55, 8'd142, 8'd108, 8'd67, 8'd132, 8'd133, 8'd81, 8'd114, 8'd66, 8'd126, 8'd153, 8'd185, 8'd212, 8'd181, 8'd152, 8'd118, 8'd90, 8'd119, 8'd160, 8'd155, 8'd143, 8'd153, 8'd141, 8'd66, 8'd131, 8'd119, 8'd56, 8'd123, 8'd69, 8'd85, 8'd149, 8'd83, 8'd123, 8'd128, 8'd157, 8'd116, 8'd99, 8'd99, 8'd135, 8'd114, 8'd153, 8'd90, 8'd161, 8'd125, 8'd124, 8'd109, 8'd111, 8'd178, 8'd144, 8'd160, 8'd117, 8'd118, 8'd137, 8'd89, 8'd95, 8'd136, 8'd173, 8'd160, 8'd134, 8'd179, 8'd139, 8'd165, 8'd153, 8'd131, 8'd122, 8'd91, 8'd134, 8'd127, 8'd149, 8'd111, 8'd160, 8'd114, 8'd167, 8'd167, 8'd188, 8'd87, 8'd99, 8'd101, 8'd180, 8'd93, 8'd151, 8'd103, 8'd96, 8'd111, 8'd122, 8'd182, 8'd175, 8'd103, 8'd112, 8'd145, 8'd78, 8'd145, 8'd132, 8'd73, 8'd124, 8'd185, 8'd174, 8'd122, 8'd77, 8'd126, 8'd84, 8'd133, 8'd129, 8'd99, 8'd130, 8'd101, 8'd190, 8'd165, 8'd171, 8'd168, 8'd80, 8'd119, 8'd112, 8'd138, 8'd166, 8'd178, 8'd91, 8'd122, 8'd79, 8'd102, 8'd117, 8'd153, 8'd113, 8'd111, 8'd131, 8'd145, 8'd53, 8'd52, 8'd86, 8'd137, 8'd123, 8'd110, 8'd164, 8'd191, 8'd111, 8'd113, 8'd186, 8'd158, 8'd157, 8'd181, 8'd153, 8'd142, 8'd163, 8'd148, 8'd152, 8'd151, 8'd140, 8'd128, 8'd136, 8'd150, 8'd123, 8'd132, 8'd152, 8'd106, 8'd127, 8'd51, 8'd77, 8'd131, 8'd78, 8'd120, 8'd93, 8'd124, 8'd175, 8'd167, 8'd137, 8'd110, 8'd185, 8'd143, 8'd120, 8'd101, 8'd182, 8'd101, 8'd146, 8'd181, 8'd131, 8'd110, 8'd83, 8'd80, 8'd133, 8'd161, 8'd128, 8'd78, 8'd81, 8'd62, 8'd32, 8'd94, 8'd75, 8'd59, 8'd76, 8'd81, 8'd164, 8'd138, 8'd112, 8'd158, 8'd113, 8'd136, 8'd113, 8'd138, 8'd184, 8'd105, 8'd131, 8'd112, 8'd104, 8'd91, 8'd135, 8'd166, 8'd148, 8'd115, 8'd105, 8'd136, 8'd38, 8'd80, 8'd85, 8'd72, 8'd92, 8'd144, 8'd132, 8'd120, 8'd118, 8'd134, 8'd114, 8'd123, 8'd159, 8'd151, 8'd93, 8'd136, 8'd87, 8'd153, 8'd77, 8'd159, 8'd135, 8'd116, 8'd75, 8'd73, 8'd107, 8'd141, 8'd90, 8'd110, 8'd120, 8'd66, 8'd121, 8'd54, 8'd69, 8'd114, 8'd126, 8'd96, 8'd95, 8'd114, 8'd118, 8'd123, 8'd138, 8'd123, 8'd120, 8'd116, 8'd113, 8'd150, 8'd132, 8'd65, 8'd70, 8'd131, 8'd155, 8'd111, 8'd106, 8'd96, 8'd130, 8'd131, 8'd128, 8'd151, 8'd64, 8'd64, 8'd124, 8'd108, 8'd70, 8'd82, 8'd148, 8'd111, 8'd58, 8'd43, 8'd69, 8'd139, 8'd89, 8'd106, 8'd142, 8'd141, 8'd87, 8'd102, 8'd129, 8'd117, 8'd168, 8'd168, 8'd150, 8'd116, 8'd82, 8'd105, 8'd150, 8'd146, 8'd101, 8'd135, 8'd140, 8'd78, 8'd121, 8'd98, 8'd140, 8'd87, 8'd141, 8'd69, 8'd158, 8'd97, 8'd80, 8'd93, 8'd137, 8'd77, 8'd160, 8'd150, 8'd139, 8'd92, 8'd97, 8'd156})
) cell_0_70 (
    .clk(clk),
    .input_index(index_0_69_70),
    .input_value(value_0_69_70),
    .input_result(result_0_69_70),
    .input_enable(enable_0_69_70),
    .output_index(index_0_70_71),
    .output_value(value_0_70_71),
    .output_result(result_0_70_71),
    .output_enable(enable_0_70_71)
);

wire [10-1:0] index_0_71_72;
wire [`DATA_WIDTH-1:0] value_0_71_72;
wire [`DATA_WIDTH*4:0] result_0_71_72;
wire enable_0_71_72;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd136, 8'd132, 8'd93, 8'd103, 8'd125, 8'd146, 8'd90, 8'd110, 8'd114, 8'd163, 8'd121, 8'd157, 8'd93, 8'd159, 8'd167, 8'd100, 8'd144, 8'd138, 8'd115, 8'd86, 8'd89, 8'd73, 8'd158, 8'd83, 8'd73, 8'd88, 8'd160, 8'd89, 8'd140, 8'd96, 8'd167, 8'd114, 8'd140, 8'd169, 8'd120, 8'd72, 8'd163, 8'd92, 8'd104, 8'd123, 8'd161, 8'd117, 8'd74, 8'd141, 8'd89, 8'd69, 8'd152, 8'd130, 8'd154, 8'd112, 8'd121, 8'd125, 8'd90, 8'd143, 8'd73, 8'd136, 8'd96, 8'd95, 8'd146, 8'd89, 8'd105, 8'd159, 8'd149, 8'd124, 8'd154, 8'd85, 8'd162, 8'd79, 8'd79, 8'd80, 8'd116, 8'd157, 8'd115, 8'd129, 8'd138, 8'd160, 8'd99, 8'd79, 8'd150, 8'd102, 8'd176, 8'd119, 8'd94, 8'd106, 8'd98, 8'd174, 8'd104, 8'd132, 8'd56, 8'd94, 8'd156, 8'd59, 8'd73, 8'd132, 8'd89, 8'd110, 8'd132, 8'd75, 8'd76, 8'd102, 8'd113, 8'd140, 8'd85, 8'd75, 8'd149, 8'd189, 8'd174, 8'd110, 8'd100, 8'd93, 8'd138, 8'd161, 8'd76, 8'd166, 8'd112, 8'd72, 8'd119, 8'd74, 8'd151, 8'd146, 8'd72, 8'd109, 8'd84, 8'd123, 8'd151, 8'd117, 8'd51, 8'd123, 8'd58, 8'd68, 8'd142, 8'd155, 8'd117, 8'd134, 8'd179, 8'd194, 8'd178, 8'd147, 8'd149, 8'd117, 8'd107, 8'd140, 8'd123, 8'd153, 8'd102, 8'd133, 8'd129, 8'd95, 8'd143, 8'd160, 8'd107, 8'd161, 8'd136, 8'd67, 8'd116, 8'd66, 8'd80, 8'd93, 8'd96, 8'd160, 8'd105, 8'd126, 8'd168, 8'd183, 8'd115, 8'd160, 8'd113, 8'd128, 8'd133, 8'd74, 8'd118, 8'd75, 8'd107, 8'd113, 8'd76, 8'd71, 8'd168, 8'd119, 8'd101, 8'd115, 8'd137, 8'd81, 8'd150, 8'd133, 8'd151, 8'd108, 8'd143, 8'd84, 8'd120, 8'd98, 8'd72, 8'd114, 8'd146, 8'd146, 8'd90, 8'd153, 8'd155, 8'd174, 8'd113, 8'd75, 8'd72, 8'd97, 8'd74, 8'd109, 8'd98, 8'd79, 8'd161, 8'd146, 8'd89, 8'd101, 8'd82, 8'd137, 8'd94, 8'd126, 8'd164, 8'd130, 8'd135, 8'd66, 8'd144, 8'd97, 8'd115, 8'd130, 8'd120, 8'd99, 8'd115, 8'd77, 8'd90, 8'd151, 8'd96, 8'd126, 8'd126, 8'd162, 8'd135, 8'd135, 8'd138, 8'd134, 8'd132, 8'd130, 8'd159, 8'd140, 8'd124, 8'd122, 8'd105, 8'd148, 8'd59, 8'd79, 8'd101, 8'd142, 8'd117, 8'd110, 8'd169, 8'd173, 8'd90, 8'd125, 8'd98, 8'd96, 8'd99, 8'd104, 8'd81, 8'd131, 8'd85, 8'd150, 8'd151, 8'd90, 8'd137, 8'd172, 8'd177, 8'd126, 8'd114, 8'd52, 8'd105, 8'd138, 8'd110, 8'd129, 8'd68, 8'd117, 8'd152, 8'd92, 8'd138, 8'd151, 8'd74, 8'd164, 8'd121, 8'd73, 8'd87, 8'd139, 8'd137, 8'd77, 8'd81, 8'd75, 8'd82, 8'd155, 8'd164, 8'd181, 8'd125, 8'd151, 8'd86, 8'd76, 8'd84, 8'd101, 8'd143, 8'd158, 8'd126, 8'd132, 8'd157, 8'd122, 8'd180, 8'd123, 8'd74, 8'd106, 8'd85, 8'd91, 8'd83, 8'd168, 8'd118, 8'd75, 8'd114, 8'd151, 8'd156, 8'd113, 8'd139, 8'd105, 8'd166, 8'd118, 8'd120, 8'd135, 8'd102, 8'd59, 8'd108, 8'd96, 8'd81, 8'd134, 8'd96, 8'd115, 8'd144, 8'd109, 8'd143, 8'd107, 8'd96, 8'd134, 8'd141, 8'd119, 8'd137, 8'd131, 8'd155, 8'd160, 8'd122, 8'd100, 8'd123, 8'd103, 8'd162, 8'd94, 8'd127, 8'd76, 8'd135, 8'd95, 8'd67, 8'd74, 8'd140, 8'd92, 8'd156, 8'd190, 8'd90, 8'd123, 8'd144, 8'd77, 8'd110, 8'd87, 8'd143, 8'd145, 8'd115, 8'd74, 8'd96, 8'd89, 8'd83, 8'd77, 8'd103, 8'd112, 8'd134, 8'd141, 8'd70, 8'd53, 8'd84, 8'd95, 8'd117, 8'd150, 8'd78, 8'd117, 8'd102, 8'd116, 8'd176, 8'd168, 8'd148, 8'd100, 8'd71, 8'd126, 8'd115, 8'd99, 8'd57, 8'd139, 8'd84, 8'd138, 8'd133, 8'd102, 8'd191, 8'd125, 8'd149, 8'd107, 8'd118, 8'd142, 8'd99, 8'd97, 8'd163, 8'd104, 8'd91, 8'd159, 8'd180, 8'd159, 8'd131, 8'd126, 8'd168, 8'd144, 8'd108, 8'd76, 8'd108, 8'd42, 8'd58, 8'd88, 8'd135, 8'd127, 8'd138, 8'd136, 8'd157, 8'd179, 8'd131, 8'd81, 8'd133, 8'd136, 8'd116, 8'd95, 8'd131, 8'd116, 8'd137, 8'd86, 8'd97, 8'd135, 8'd156, 8'd147, 8'd92, 8'd127, 8'd103, 8'd71, 8'd121, 8'd56, 8'd98, 8'd76, 8'd59, 8'd120, 8'd122, 8'd130, 8'd165, 8'd118, 8'd134, 8'd74, 8'd146, 8'd129, 8'd73, 8'd89, 8'd116, 8'd133, 8'd160, 8'd164, 8'd121, 8'd103, 8'd109, 8'd114, 8'd101, 8'd121, 8'd117, 8'd72, 8'd98, 8'd123, 8'd155, 8'd150, 8'd60, 8'd88, 8'd77, 8'd164, 8'd199, 8'd143, 8'd109, 8'd126, 8'd125, 8'd90, 8'd97, 8'd81, 8'd145, 8'd69, 8'd72, 8'd88, 8'd101, 8'd144, 8'd95, 8'd104, 8'd123, 8'd165, 8'd108, 8'd125, 8'd146, 8'd152, 8'd157, 8'd80, 8'd152, 8'd96, 8'd170, 8'd168, 8'd128, 8'd78, 8'd101, 8'd76, 8'd150, 8'd155, 8'd120, 8'd100, 8'd158, 8'd137, 8'd152, 8'd132, 8'd149, 8'd184, 8'd124, 8'd116, 8'd134, 8'd112, 8'd131, 8'd141, 8'd65, 8'd100, 8'd103, 8'd107, 8'd104, 8'd110, 8'd155, 8'd87, 8'd133, 8'd152, 8'd74, 8'd135, 8'd101, 8'd92, 8'd157, 8'd147, 8'd152, 8'd105, 8'd137, 8'd103, 8'd106, 8'd168, 8'd146, 8'd133, 8'd127, 8'd112, 8'd102, 8'd98, 8'd140, 8'd87, 8'd162, 8'd83, 8'd158, 8'd128, 8'd102, 8'd75, 8'd124, 8'd78, 8'd68, 8'd112, 8'd149, 8'd127, 8'd97, 8'd140, 8'd77, 8'd158, 8'd157, 8'd145, 8'd126, 8'd114, 8'd168, 8'd103, 8'd101, 8'd135, 8'd97, 8'd171, 8'd171, 8'd125, 8'd98, 8'd70, 8'd136, 8'd124, 8'd121, 8'd74, 8'd93, 8'd49, 8'd57, 8'd91, 8'd125, 8'd120, 8'd85, 8'd135, 8'd138, 8'd115, 8'd187, 8'd108, 8'd169, 8'd93, 8'd132, 8'd124, 8'd85, 8'd90, 8'd107, 8'd105, 8'd126, 8'd144, 8'd188, 8'd110, 8'd159, 8'd129, 8'd145, 8'd148, 8'd73, 8'd90, 8'd132, 8'd69, 8'd98, 8'd124, 8'd107, 8'd153, 8'd96, 8'd140, 8'd108, 8'd189, 8'd89, 8'd106, 8'd119, 8'd86, 8'd130, 8'd94, 8'd165, 8'd182, 8'd148, 8'd158, 8'd164, 8'd152, 8'd169, 8'd94, 8'd107, 8'd122, 8'd104, 8'd141, 8'd134, 8'd169, 8'd121, 8'd139, 8'd162, 8'd167, 8'd90, 8'd129, 8'd129, 8'd94, 8'd167, 8'd112, 8'd132, 8'd161, 8'd121, 8'd109, 8'd138, 8'd61, 8'd63, 8'd157, 8'd171, 8'd182, 8'd163, 8'd101, 8'd190, 8'd154, 8'd161, 8'd186, 8'd97, 8'd124, 8'd100, 8'd94, 8'd81, 8'd116, 8'd94, 8'd160, 8'd143, 8'd88, 8'd112, 8'd104, 8'd123, 8'd101, 8'd161, 8'd77, 8'd167, 8'd72, 8'd101, 8'd96, 8'd70, 8'd110, 8'd184, 8'd119, 8'd143, 8'd135, 8'd128, 8'd112, 8'd100, 8'd80, 8'd83, 8'd46, 8'd106, 8'd45, 8'd135, 8'd96, 8'd142, 8'd125, 8'd112, 8'd115, 8'd120, 8'd101, 8'd97, 8'd110, 8'd130, 8'd138, 8'd81, 8'd112, 8'd149, 8'd125, 8'd148, 8'd111, 8'd78, 8'd143, 8'd158, 8'd115, 8'd63, 8'd73, 8'd127, 8'd72, 8'd80, 8'd134, 8'd127, 8'd95, 8'd141, 8'd159, 8'd87, 8'd104, 8'd89, 8'd78, 8'd155, 8'd106, 8'd89, 8'd161, 8'd144, 8'd124, 8'd144, 8'd105, 8'd139, 8'd152, 8'd140, 8'd166, 8'd87, 8'd110, 8'd126, 8'd76, 8'd153, 8'd137, 8'd87, 8'd104, 8'd162, 8'd164, 8'd130, 8'd164, 8'd137, 8'd101, 8'd163, 8'd116})
) cell_0_71 (
    .clk(clk),
    .input_index(index_0_70_71),
    .input_value(value_0_70_71),
    .input_result(result_0_70_71),
    .input_enable(enable_0_70_71),
    .output_index(index_0_71_72),
    .output_value(value_0_71_72),
    .output_result(result_0_71_72),
    .output_enable(enable_0_71_72)
);

wire [10-1:0] index_0_72_73;
wire [`DATA_WIDTH-1:0] value_0_72_73;
wire [`DATA_WIDTH*4:0] result_0_72_73;
wire enable_0_72_73;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd102, 8'd154, 8'd89, 8'd119, 8'd134, 8'd77, 8'd144, 8'd107, 8'd85, 8'd65, 8'd89, 8'd114, 8'd115, 8'd83, 8'd126, 8'd82, 8'd58, 8'd68, 8'd78, 8'd122, 8'd151, 8'd133, 8'd105, 8'd115, 8'd81, 8'd164, 8'd104, 8'd124, 8'd73, 8'd132, 8'd145, 8'd116, 8'd148, 8'd93, 8'd105, 8'd115, 8'd106, 8'd97, 8'd95, 8'd4, 8'd45, 8'd55, 8'd16, 8'd81, 8'd27, 8'd84, 8'd62, 8'd95, 8'd64, 8'd94, 8'd128, 8'd121, 8'd75, 8'd163, 8'd145, 8'd76, 8'd118, 8'd109, 8'd146, 8'd55, 8'd56, 8'd124, 8'd71, 8'd102, 8'd91, 8'd42, 8'd34, 8'd67, 8'd43, 8'd80, 8'd98, 8'd101, 8'd84, 8'd135, 8'd75, 8'd65, 8'd48, 8'd83, 8'd51, 8'd88, 8'd103, 8'd161, 8'd81, 8'd153, 8'd91, 8'd78, 8'd99, 8'd175, 8'd154, 8'd133, 8'd108, 8'd130, 8'd80, 8'd93, 8'd74, 8'd129, 8'd162, 8'd90, 8'd112, 8'd148, 8'd147, 8'd78, 8'd82, 8'd87, 8'd107, 8'd70, 8'd107, 8'd126, 8'd148, 8'd130, 8'd159, 8'd138, 8'd122, 8'd132, 8'd86, 8'd100, 8'd97, 8'd130, 8'd144, 8'd116, 8'd119, 8'd150, 8'd147, 8'd156, 8'd123, 8'd101, 8'd103, 8'd75, 8'd91, 8'd109, 8'd166, 8'd159, 8'd180, 8'd84, 8'd68, 8'd155, 8'd134, 8'd100, 8'd123, 8'd143, 8'd86, 8'd100, 8'd127, 8'd94, 8'd93, 8'd172, 8'd106, 8'd128, 8'd115, 8'd164, 8'd115, 8'd89, 8'd91, 8'd84, 8'd155, 8'd102, 8'd85, 8'd170, 8'd134, 8'd87, 8'd152, 8'd107, 8'd137, 8'd166, 8'd97, 8'd135, 8'd152, 8'd138, 8'd138, 8'd127, 8'd85, 8'd180, 8'd98, 8'd138, 8'd143, 8'd120, 8'd105, 8'd114, 8'd109, 8'd128, 8'd96, 8'd134, 8'd71, 8'd92, 8'd160, 8'd146, 8'd91, 8'd92, 8'd166, 8'd91, 8'd172, 8'd88, 8'd181, 8'd89, 8'd109, 8'd161, 8'd136, 8'd144, 8'd130, 8'd102, 8'd167, 8'd155, 8'd153, 8'd128, 8'd143, 8'd134, 8'd71, 8'd113, 8'd130, 8'd72, 8'd139, 8'd136, 8'd117, 8'd71, 8'd127, 8'd109, 8'd168, 8'd169, 8'd146, 8'd113, 8'd160, 8'd122, 8'd118, 8'd119, 8'd114, 8'd106, 8'd190, 8'd119, 8'd75, 8'd141, 8'd121, 8'd134, 8'd140, 8'd107, 8'd141, 8'd151, 8'd152, 8'd103, 8'd130, 8'd122, 8'd66, 8'd119, 8'd136, 8'd92, 8'd90, 8'd110, 8'd117, 8'd129, 8'd100, 8'd119, 8'd100, 8'd119, 8'd138, 8'd106, 8'd150, 8'd160, 8'd127, 8'd83, 8'd149, 8'd109, 8'd94, 8'd97, 8'd129, 8'd162, 8'd123, 8'd185, 8'd117, 8'd165, 8'd162, 8'd103, 8'd130, 8'd169, 8'd139, 8'd122, 8'd152, 8'd149, 8'd81, 8'd100, 8'd84, 8'd87, 8'd156, 8'd131, 8'd174, 8'd150, 8'd74, 8'd122, 8'd148, 8'd132, 8'd89, 8'd86, 8'd106, 8'd135, 8'd134, 8'd158, 8'd106, 8'd154, 8'd144, 8'd164, 8'd111, 8'd131, 8'd127, 8'd154, 8'd110, 8'd131, 8'd152, 8'd73, 8'd98, 8'd128, 8'd103, 8'd201, 8'd130, 8'd97, 8'd115, 8'd144, 8'd145, 8'd116, 8'd117, 8'd142, 8'd158, 8'd150, 8'd123, 8'd181, 8'd90, 8'd139, 8'd81, 8'd159, 8'd162, 8'd143, 8'd161, 8'd171, 8'd176, 8'd126, 8'd152, 8'd72, 8'd138, 8'd165, 8'd139, 8'd199, 8'd143, 8'd144, 8'd142, 8'd97, 8'd89, 8'd75, 8'd109, 8'd147, 8'd116, 8'd167, 8'd116, 8'd127, 8'd99, 8'd125, 8'd70, 8'd92, 8'd117, 8'd96, 8'd103, 8'd121, 8'd90, 8'd95, 8'd123, 8'd132, 8'd160, 8'd143, 8'd116, 8'd204, 8'd191, 8'd81, 8'd104, 8'd105, 8'd157, 8'd99, 8'd174, 8'd120, 8'd160, 8'd93, 8'd130, 8'd121, 8'd167, 8'd153, 8'd84, 8'd118, 8'd95, 8'd87, 8'd169, 8'd91, 8'd126, 8'd143, 8'd131, 8'd100, 8'd135, 8'd121, 8'd101, 8'd195, 8'd158, 8'd120, 8'd105, 8'd99, 8'd167, 8'd148, 8'd88, 8'd108, 8'd122, 8'd88, 8'd125, 8'd163, 8'd126, 8'd110, 8'd139, 8'd109, 8'd122, 8'd154, 8'd83, 8'd125, 8'd118, 8'd69, 8'd64, 8'd101, 8'd117, 8'd82, 8'd89, 8'd145, 8'd107, 8'd113, 8'd153, 8'd170, 8'd113, 8'd164, 8'd179, 8'd124, 8'd134, 8'd111, 8'd107, 8'd128, 8'd82, 8'd67, 8'd109, 8'd158, 8'd87, 8'd128, 8'd139, 8'd120, 8'd128, 8'd61, 8'd112, 8'd58, 8'd97, 8'd97, 8'd130, 8'd69, 8'd123, 8'd85, 8'd146, 8'd88, 8'd160, 8'd159, 8'd119, 8'd101, 8'd105, 8'd121, 8'd93, 8'd64, 8'd115, 8'd54, 8'd148, 8'd101, 8'd70, 8'd142, 8'd85, 8'd137, 8'd151, 8'd62, 8'd115, 8'd102, 8'd57, 8'd83, 8'd157, 8'd111, 8'd59, 8'd113, 8'd87, 8'd72, 8'd115, 8'd143, 8'd178, 8'd149, 8'd175, 8'd105, 8'd134, 8'd99, 8'd67, 8'd133, 8'd141, 8'd58, 8'd67, 8'd82, 8'd118, 8'd77, 8'd87, 8'd91, 8'd126, 8'd144, 8'd146, 8'd124, 8'd62, 8'd112, 8'd106, 8'd67, 8'd122, 8'd125, 8'd130, 8'd91, 8'd154, 8'd190, 8'd140, 8'd173, 8'd79, 8'd94, 8'd94, 8'd129, 8'd100, 8'd162, 8'd86, 8'd86, 8'd87, 8'd92, 8'd175, 8'd168, 8'd118, 8'd81, 8'd59, 8'd101, 8'd95, 8'd147, 8'd51, 8'd96, 8'd146, 8'd136, 8'd79, 8'd138, 8'd106, 8'd121, 8'd89, 8'd108, 8'd129, 8'd83, 8'd80, 8'd80, 8'd136, 8'd114, 8'd99, 8'd101, 8'd95, 8'd88, 8'd97, 8'd105, 8'd124, 8'd81, 8'd76, 8'd123, 8'd144, 8'd125, 8'd95, 8'd54, 8'd156, 8'd131, 8'd83, 8'd140, 8'd112, 8'd159, 8'd67, 8'd120, 8'd91, 8'd108, 8'd101, 8'd80, 8'd111, 8'd73, 8'd74, 8'd100, 8'd112, 8'd112, 8'd105, 8'd156, 8'd168, 8'd83, 8'd170, 8'd125, 8'd128, 8'd100, 8'd59, 8'd89, 8'd99, 8'd148, 8'd157, 8'd83, 8'd127, 8'd94, 8'd113, 8'd155, 8'd77, 8'd69, 8'd131, 8'd139, 8'd153, 8'd99, 8'd140, 8'd162, 8'd157, 8'd145, 8'd162, 8'd176, 8'd177, 8'd138, 8'd169, 8'd156, 8'd156, 8'd50, 8'd73, 8'd142, 8'd80, 8'd130, 8'd120, 8'd161, 8'd128, 8'd174, 8'd96, 8'd132, 8'd135, 8'd107, 8'd169, 8'd153, 8'd147, 8'd93, 8'd84, 8'd139, 8'd114, 8'd117, 8'd128, 8'd167, 8'd146, 8'd89, 8'd113, 8'd95, 8'd65, 8'd128, 8'd106, 8'd70, 8'd54, 8'd82, 8'd97, 8'd65, 8'd54, 8'd108, 8'd90, 8'd144, 8'd154, 8'd159, 8'd112, 8'd158, 8'd148, 8'd99, 8'd89, 8'd160, 8'd83, 8'd164, 8'd149, 8'd163, 8'd138, 8'd74, 8'd152, 8'd156, 8'd85, 8'd89, 8'd156, 8'd97, 8'd43, 8'd30, 8'd61, 8'd78, 8'd115, 8'd87, 8'd97, 8'd107, 8'd121, 8'd118, 8'd71, 8'd94, 8'd165, 8'd74, 8'd88, 8'd136, 8'd156, 8'd145, 8'd88, 8'd146, 8'd74, 8'd101, 8'd153, 8'd83, 8'd71, 8'd131, 8'd128, 8'd108, 8'd76, 8'd103, 8'd72, 8'd121, 8'd85, 8'd139, 8'd124, 8'd114, 8'd98, 8'd67, 8'd111, 8'd144, 8'd107, 8'd132, 8'd144, 8'd81, 8'd131, 8'd104, 8'd79, 8'd140, 8'd81, 8'd89, 8'd153, 8'd93, 8'd111, 8'd85, 8'd117, 8'd123, 8'd73, 8'd142, 8'd63, 8'd80, 8'd136, 8'd49, 8'd124, 8'd160, 8'd150, 8'd161, 8'd75, 8'd104, 8'd64, 8'd91, 8'd133, 8'd147, 8'd117, 8'd146, 8'd139, 8'd100, 8'd86, 8'd145, 8'd86, 8'd155, 8'd70, 8'd97, 8'd169, 8'd96, 8'd137, 8'd125, 8'd78, 8'd124, 8'd87, 8'd167, 8'd154, 8'd147, 8'd80, 8'd138, 8'd136, 8'd149, 8'd159, 8'd92, 8'd114, 8'd166, 8'd166, 8'd90, 8'd162, 8'd73, 8'd143, 8'd119, 8'd70, 8'd125})
) cell_0_72 (
    .clk(clk),
    .input_index(index_0_71_72),
    .input_value(value_0_71_72),
    .input_result(result_0_71_72),
    .input_enable(enable_0_71_72),
    .output_index(index_0_72_73),
    .output_value(value_0_72_73),
    .output_result(result_0_72_73),
    .output_enable(enable_0_72_73)
);

wire [10-1:0] index_0_73_74;
wire [`DATA_WIDTH-1:0] value_0_73_74;
wire [`DATA_WIDTH*4:0] result_0_73_74;
wire enable_0_73_74;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd141, 8'd163, 8'd109, 8'd102, 8'd79, 8'd149, 8'd107, 8'd61, 8'd103, 8'd110, 8'd114, 8'd133, 8'd112, 8'd85, 8'd88, 8'd114, 8'd88, 8'd68, 8'd89, 8'd108, 8'd72, 8'd72, 8'd86, 8'd146, 8'd106, 8'd167, 8'd128, 8'd95, 8'd163, 8'd136, 8'd72, 8'd153, 8'd68, 8'd113, 8'd103, 8'd60, 8'd135, 8'd57, 8'd132, 8'd110, 8'd78, 8'd100, 8'd50, 8'd69, 8'd69, 8'd51, 8'd101, 8'd113, 8'd107, 8'd130, 8'd134, 8'd71, 8'd112, 8'd118, 8'd76, 8'd158, 8'd117, 8'd156, 8'd156, 8'd154, 8'd170, 8'd135, 8'd132, 8'd50, 8'd81, 8'd120, 8'd140, 8'd150, 8'd116, 8'd128, 8'd137, 8'd101, 8'd68, 8'd102, 8'd50, 8'd34, 8'd55, 8'd123, 8'd112, 8'd64, 8'd86, 8'd127, 8'd125, 8'd142, 8'd100, 8'd86, 8'd112, 8'd138, 8'd112, 8'd120, 8'd135, 8'd68, 8'd131, 8'd104, 8'd155, 8'd155, 8'd88, 8'd138, 8'd73, 8'd119, 8'd112, 8'd132, 8'd93, 8'd117, 8'd91, 8'd93, 8'd65, 8'd65, 8'd120, 8'd110, 8'd80, 8'd105, 8'd99, 8'd124, 8'd155, 8'd156, 8'd97, 8'd153, 8'd147, 8'd117, 8'd99, 8'd101, 8'd134, 8'd161, 8'd116, 8'd144, 8'd108, 8'd148, 8'd149, 8'd150, 8'd141, 8'd149, 8'd105, 8'd84, 8'd106, 8'd97, 8'd151, 8'd89, 8'd97, 8'd141, 8'd84, 8'd175, 8'd178, 8'd118, 8'd92, 8'd102, 8'd119, 8'd135, 8'd173, 8'd119, 8'd133, 8'd173, 8'd153, 8'd125, 8'd109, 8'd102, 8'd180, 8'd161, 8'd155, 8'd175, 8'd184, 8'd141, 8'd140, 8'd139, 8'd115, 8'd113, 8'd163, 8'd139, 8'd108, 8'd159, 8'd100, 8'd135, 8'd133, 8'd195, 8'd97, 8'd130, 8'd143, 8'd96, 8'd168, 8'd110, 8'd118, 8'd94, 8'd103, 8'd88, 8'd113, 8'd164, 8'd152, 8'd150, 8'd145, 8'd190, 8'd182, 8'd150, 8'd188, 8'd85, 8'd88, 8'd128, 8'd119, 8'd105, 8'd93, 8'd177, 8'd172, 8'd150, 8'd176, 8'd116, 8'd131, 8'd153, 8'd102, 8'd83, 8'd113, 8'd111, 8'd99, 8'd129, 8'd181, 8'd119, 8'd161, 8'd168, 8'd145, 8'd174, 8'd117, 8'd142, 8'd177, 8'd115, 8'd161, 8'd96, 8'd165, 8'd149, 8'd190, 8'd134, 8'd158, 8'd145, 8'd130, 8'd139, 8'd147, 8'd111, 8'd133, 8'd104, 8'd84, 8'd96, 8'd182, 8'd157, 8'd172, 8'd108, 8'd184, 8'd150, 8'd112, 8'd107, 8'd202, 8'd173, 8'd141, 8'd122, 8'd107, 8'd171, 8'd90, 8'd111, 8'd132, 8'd132, 8'd185, 8'd185, 8'd122, 8'd146, 8'd99, 8'd74, 8'd79, 8'd156, 8'd97, 8'd170, 8'd131, 8'd102, 8'd139, 8'd101, 8'd112, 8'd136, 8'd93, 8'd198, 8'd187, 8'd204, 8'd189, 8'd174, 8'd145, 8'd149, 8'd97, 8'd196, 8'd150, 8'd130, 8'd125, 8'd160, 8'd114, 8'd119, 8'd106, 8'd128, 8'd114, 8'd82, 8'd106, 8'd135, 8'd163, 8'd150, 8'd109, 8'd102, 8'd64, 8'd54, 8'd149, 8'd141, 8'd132, 8'd198, 8'd155, 8'd130, 8'd154, 8'd105, 8'd178, 8'd147, 8'd178, 8'd122, 8'd104, 8'd108, 8'd145, 8'd111, 8'd142, 8'd87, 8'd104, 8'd56, 8'd66, 8'd123, 8'd142, 8'd146, 8'd65, 8'd125, 8'd119, 8'd130, 8'd87, 8'd90, 8'd67, 8'd141, 8'd159, 8'd101, 8'd79, 8'd69, 8'd165, 8'd164, 8'd166, 8'd90, 8'd159, 8'd96, 8'd50, 8'd67, 8'd48, 8'd97, 8'd73, 8'd108, 8'd118, 8'd159, 8'd130, 8'd167, 8'd71, 8'd84, 8'd138, 8'd88, 8'd134, 8'd117, 8'd108, 8'd93, 8'd128, 8'd124, 8'd130, 8'd96, 8'd125, 8'd132, 8'd157, 8'd118, 8'd55, 8'd45, 8'd80, 8'd114, 8'd123, 8'd75, 8'd74, 8'd54, 8'd89, 8'd154, 8'd146, 8'd112, 8'd133, 8'd71, 8'd79, 8'd131, 8'd109, 8'd49, 8'd120, 8'd100, 8'd63, 8'd165, 8'd120, 8'd140, 8'd124, 8'd151, 8'd147, 8'd121, 8'd122, 8'd26, 8'd33, 8'd54, 8'd69, 8'd117, 8'd60, 8'd62, 8'd101, 8'd127, 8'd200, 8'd173, 8'd116, 8'd102, 8'd50, 8'd140, 8'd80, 8'd109, 8'd106, 8'd83, 8'd120, 8'd72, 8'd159, 8'd172, 8'd170, 8'd180, 8'd105, 8'd61, 8'd125, 8'd61, 8'd72, 8'd43, 8'd62, 8'd87, 8'd107, 8'd70, 8'd107, 8'd113, 8'd126, 8'd161, 8'd86, 8'd76, 8'd78, 8'd65, 8'd66, 8'd96, 8'd149, 8'd66, 8'd151, 8'd74, 8'd134, 8'd154, 8'd144, 8'd132, 8'd206, 8'd149, 8'd107, 8'd138, 8'd106, 8'd75, 8'd46, 8'd56, 8'd126, 8'd98, 8'd132, 8'd174, 8'd126, 8'd125, 8'd108, 8'd117, 8'd143, 8'd72, 8'd135, 8'd117, 8'd84, 8'd149, 8'd121, 8'd140, 8'd103, 8'd89, 8'd105, 8'd208, 8'd177, 8'd149, 8'd181, 8'd138, 8'd140, 8'd147, 8'd109, 8'd143, 8'd117, 8'd114, 8'd151, 8'd151, 8'd96, 8'd96, 8'd108, 8'd147, 8'd146, 8'd111, 8'd98, 8'd108, 8'd126, 8'd126, 8'd152, 8'd122, 8'd129, 8'd69, 8'd139, 8'd182, 8'd242, 8'd233, 8'd172, 8'd169, 8'd158, 8'd152, 8'd115, 8'd152, 8'd94, 8'd84, 8'd107, 8'd108, 8'd101, 8'd76, 8'd125, 8'd101, 8'd96, 8'd130, 8'd81, 8'd115, 8'd173, 8'd178, 8'd125, 8'd124, 8'd76, 8'd148, 8'd179, 8'd142, 8'd162, 8'd144, 8'd197, 8'd178, 8'd132, 8'd120, 8'd170, 8'd109, 8'd88, 8'd157, 8'd123, 8'd124, 8'd71, 8'd159, 8'd152, 8'd134, 8'd135, 8'd118, 8'd94, 8'd99, 8'd94, 8'd99, 8'd123, 8'd137, 8'd85, 8'd108, 8'd79, 8'd96, 8'd132, 8'd175, 8'd193, 8'd110, 8'd143, 8'd91, 8'd136, 8'd125, 8'd78, 8'd80, 8'd75, 8'd80, 8'd123, 8'd124, 8'd128, 8'd79, 8'd128, 8'd85, 8'd89, 8'd101, 8'd97, 8'd131, 8'd130, 8'd139, 8'd152, 8'd77, 8'd122, 8'd102, 8'd169, 8'd140, 8'd121, 8'd121, 8'd116, 8'd116, 8'd136, 8'd159, 8'd129, 8'd129, 8'd81, 8'd149, 8'd99, 8'd86, 8'd118, 8'd66, 8'd76, 8'd108, 8'd70, 8'd136, 8'd142, 8'd84, 8'd158, 8'd97, 8'd118, 8'd77, 8'd155, 8'd160, 8'd106, 8'd141, 8'd106, 8'd158, 8'd112, 8'd193, 8'd167, 8'd159, 8'd183, 8'd190, 8'd127, 8'd144, 8'd122, 8'd122, 8'd138, 8'd114, 8'd150, 8'd158, 8'd112, 8'd147, 8'd159, 8'd152, 8'd171, 8'd82, 8'd99, 8'd105, 8'd128, 8'd112, 8'd164, 8'd123, 8'd130, 8'd63, 8'd78, 8'd151, 8'd165, 8'd99, 8'd167, 8'd175, 8'd121, 8'd125, 8'd142, 8'd207, 8'd189, 8'd149, 8'd178, 8'd75, 8'd161, 8'd98, 8'd111, 8'd66, 8'd108, 8'd130, 8'd82, 8'd156, 8'd92, 8'd101, 8'd163, 8'd136, 8'd119, 8'd64, 8'd85, 8'd99, 8'd135, 8'd83, 8'd71, 8'd163, 8'd135, 8'd109, 8'd173, 8'd97, 8'd106, 8'd123, 8'd149, 8'd75, 8'd140, 8'd122, 8'd87, 8'd160, 8'd167, 8'd150, 8'd142, 8'd86, 8'd155, 8'd168, 8'd97, 8'd79, 8'd138, 8'd51, 8'd131, 8'd143, 8'd86, 8'd99, 8'd77, 8'd96, 8'd116, 8'd141, 8'd97, 8'd146, 8'd104, 8'd66, 8'd111, 8'd75, 8'd106, 8'd112, 8'd125, 8'd132, 8'd99, 8'd98, 8'd81, 8'd110, 8'd160, 8'd152, 8'd109, 8'd149, 8'd141, 8'd147, 8'd137, 8'd62, 8'd145, 8'd123, 8'd114, 8'd181, 8'd101, 8'd129, 8'd132, 8'd142, 8'd73, 8'd71, 8'd129, 8'd139, 8'd67, 8'd78, 8'd125, 8'd67, 8'd100, 8'd168, 8'd110, 8'd98, 8'd110, 8'd120, 8'd77, 8'd141, 8'd156, 8'd160, 8'd80, 8'd111, 8'd116, 8'd91, 8'd136, 8'd92, 8'd93, 8'd116, 8'd76, 8'd162, 8'd136, 8'd149, 8'd162, 8'd157, 8'd146, 8'd98, 8'd128, 8'd133, 8'd158, 8'd144, 8'd143, 8'd166})
) cell_0_73 (
    .clk(clk),
    .input_index(index_0_72_73),
    .input_value(value_0_72_73),
    .input_result(result_0_72_73),
    .input_enable(enable_0_72_73),
    .output_index(index_0_73_74),
    .output_value(value_0_73_74),
    .output_result(result_0_73_74),
    .output_enable(enable_0_73_74)
);

wire [10-1:0] index_0_74_75;
wire [`DATA_WIDTH-1:0] value_0_74_75;
wire [`DATA_WIDTH*4:0] result_0_74_75;
wire enable_0_74_75;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd155, 8'd162, 8'd141, 8'd119, 8'd97, 8'd129, 8'd172, 8'd115, 8'd135, 8'd174, 8'd162, 8'd133, 8'd103, 8'd179, 8'd132, 8'd176, 8'd104, 8'd107, 8'd81, 8'd140, 8'd166, 8'd137, 8'd151, 8'd106, 8'd158, 8'd147, 8'd116, 8'd117, 8'd161, 8'd126, 8'd93, 8'd163, 8'd89, 8'd96, 8'd121, 8'd77, 8'd147, 8'd156, 8'd169, 8'd128, 8'd116, 8'd100, 8'd153, 8'd94, 8'd156, 8'd145, 8'd96, 8'd111, 8'd126, 8'd77, 8'd65, 8'd93, 8'd94, 8'd80, 8'd146, 8'd146, 8'd74, 8'd138, 8'd82, 8'd80, 8'd161, 8'd101, 8'd147, 8'd123, 8'd115, 8'd161, 8'd136, 8'd125, 8'd171, 8'd109, 8'd171, 8'd179, 8'd157, 8'd112, 8'd166, 8'd101, 8'd77, 8'd121, 8'd113, 8'd105, 8'd110, 8'd74, 8'd117, 8'd93, 8'd146, 8'd163, 8'd159, 8'd90, 8'd126, 8'd85, 8'd119, 8'd97, 8'd118, 8'd98, 8'd112, 8'd186, 8'd180, 8'd135, 8'd120, 8'd188, 8'd152, 8'd93, 8'd116, 8'd161, 8'd91, 8'd135, 8'd159, 8'd140, 8'd130, 8'd115, 8'd115, 8'd129, 8'd166, 8'd135, 8'd106, 8'd90, 8'd112, 8'd150, 8'd160, 8'd144, 8'd77, 8'd89, 8'd145, 8'd163, 8'd130, 8'd170, 8'd144, 8'd131, 8'd126, 8'd111, 8'd62, 8'd56, 8'd69, 8'd144, 8'd113, 8'd175, 8'd145, 8'd57, 8'd160, 8'd87, 8'd121, 8'd129, 8'd131, 8'd152, 8'd156, 8'd67, 8'd155, 8'd74, 8'd112, 8'd161, 8'd164, 8'd119, 8'd115, 8'd149, 8'd113, 8'd165, 8'd155, 8'd97, 8'd77, 8'd115, 8'd98, 8'd110, 8'd134, 8'd78, 8'd126, 8'd58, 8'd71, 8'd135, 8'd134, 8'd125, 8'd129, 8'd151, 8'd156, 8'd134, 8'd85, 8'd164, 8'd111, 8'd78, 8'd113, 8'd133, 8'd162, 8'd109, 8'd160, 8'd105, 8'd161, 8'd99, 8'd101, 8'd70, 8'd95, 8'd63, 8'd63, 8'd125, 8'd62, 8'd104, 8'd159, 8'd87, 8'd142, 8'd125, 8'd112, 8'd104, 8'd137, 8'd164, 8'd101, 8'd133, 8'd103, 8'd75, 8'd120, 8'd154, 8'd112, 8'd97, 8'd89, 8'd185, 8'd169, 8'd74, 8'd117, 8'd64, 8'd131, 8'd75, 8'd112, 8'd101, 8'd136, 8'd160, 8'd123, 8'd125, 8'd75, 8'd108, 8'd105, 8'd139, 8'd86, 8'd87, 8'd128, 8'd77, 8'd75, 8'd102, 8'd132, 8'd92, 8'd147, 8'd153, 8'd106, 8'd177, 8'd154, 8'd85, 8'd129, 8'd80, 8'd84, 8'd152, 8'd101, 8'd52, 8'd67, 8'd100, 8'd167, 8'd89, 8'd107, 8'd145, 8'd95, 8'd131, 8'd117, 8'd111, 8'd65, 8'd136, 8'd146, 8'd168, 8'd112, 8'd155, 8'd126, 8'd201, 8'd122, 8'd206, 8'd119, 8'd117, 8'd143, 8'd77, 8'd88, 8'd131, 8'd115, 8'd131, 8'd71, 8'd117, 8'd139, 8'd151, 8'd132, 8'd98, 8'd71, 8'd107, 8'd94, 8'd119, 8'd77, 8'd114, 8'd93, 8'd154, 8'd102, 8'd177, 8'd101, 8'd183, 8'd193, 8'd150, 8'd128, 8'd87, 8'd123, 8'd108, 8'd89, 8'd59, 8'd129, 8'd139, 8'd102, 8'd134, 8'd157, 8'd121, 8'd96, 8'd130, 8'd97, 8'd118, 8'd89, 8'd147, 8'd121, 8'd140, 8'd169, 8'd174, 8'd123, 8'd97, 8'd187, 8'd210, 8'd137, 8'd169, 8'd158, 8'd140, 8'd45, 8'd54, 8'd74, 8'd99, 8'd124, 8'd95, 8'd154, 8'd111, 8'd71, 8'd132, 8'd67, 8'd155, 8'd115, 8'd64, 8'd129, 8'd140, 8'd163, 8'd125, 8'd104, 8'd97, 8'd148, 8'd128, 8'd210, 8'd218, 8'd180, 8'd140, 8'd150, 8'd132, 8'd111, 8'd106, 8'd118, 8'd156, 8'd66, 8'd159, 8'd142, 8'd168, 8'd112, 8'd137, 8'd85, 8'd79, 8'd132, 8'd104, 8'd100, 8'd122, 8'd99, 8'd167, 8'd86, 8'd131, 8'd120, 8'd134, 8'd137, 8'd131, 8'd100, 8'd79, 8'd123, 8'd121, 8'd102, 8'd89, 8'd81, 8'd148, 8'd82, 8'd169, 8'd110, 8'd106, 8'd94, 8'd141, 8'd122, 8'd81, 8'd166, 8'd135, 8'd88, 8'd99, 8'd119, 8'd123, 8'd158, 8'd93, 8'd165, 8'd140, 8'd144, 8'd125, 8'd85, 8'd162, 8'd115, 8'd126, 8'd134, 8'd125, 8'd84, 8'd160, 8'd109, 8'd89, 8'd157, 8'd120, 8'd129, 8'd150, 8'd123, 8'd141, 8'd176, 8'd92, 8'd111, 8'd75, 8'd68, 8'd144, 8'd146, 8'd90, 8'd112, 8'd195, 8'd162, 8'd125, 8'd89, 8'd122, 8'd173, 8'd159, 8'd116, 8'd155, 8'd130, 8'd172, 8'd82, 8'd103, 8'd186, 8'd150, 8'd129, 8'd145, 8'd144, 8'd171, 8'd195, 8'd85, 8'd89, 8'd146, 8'd141, 8'd147, 8'd64, 8'd116, 8'd142, 8'd146, 8'd153, 8'd161, 8'd153, 8'd135, 8'd168, 8'd175, 8'd197, 8'd168, 8'd176, 8'd165, 8'd165, 8'd106, 8'd130, 8'd118, 8'd104, 8'd104, 8'd131, 8'd208, 8'd150, 8'd141, 8'd104, 8'd125, 8'd74, 8'd88, 8'd116, 8'd101, 8'd73, 8'd123, 8'd116, 8'd105, 8'd93, 8'd186, 8'd148, 8'd196, 8'd139, 8'd144, 8'd121, 8'd172, 8'd178, 8'd126, 8'd132, 8'd126, 8'd150, 8'd108, 8'd169, 8'd169, 8'd173, 8'd162, 8'd174, 8'd97, 8'd155, 8'd105, 8'd118, 8'd72, 8'd75, 8'd78, 8'd108, 8'd63, 8'd125, 8'd96, 8'd128, 8'd135, 8'd129, 8'd159, 8'd147, 8'd91, 8'd103, 8'd107, 8'd104, 8'd176, 8'd142, 8'd166, 8'd173, 8'd194, 8'd167, 8'd147, 8'd125, 8'd153, 8'd163, 8'd84, 8'd140, 8'd129, 8'd112, 8'd102, 8'd99, 8'd137, 8'd98, 8'd93, 8'd114, 8'd108, 8'd121, 8'd143, 8'd131, 8'd176, 8'd157, 8'd181, 8'd113, 8'd126, 8'd130, 8'd84, 8'd125, 8'd127, 8'd215, 8'd148, 8'd106, 8'd124, 8'd145, 8'd75, 8'd82, 8'd56, 8'd128, 8'd65, 8'd120, 8'd67, 8'd79, 8'd89, 8'd169, 8'd180, 8'd173, 8'd169, 8'd169, 8'd120, 8'd140, 8'd123, 8'd130, 8'd131, 8'd127, 8'd159, 8'd182, 8'd187, 8'd156, 8'd167, 8'd126, 8'd149, 8'd122, 8'd137, 8'd73, 8'd64, 8'd58, 8'd75, 8'd133, 8'd88, 8'd115, 8'd156, 8'd137, 8'd112, 8'd125, 8'd138, 8'd115, 8'd144, 8'd86, 8'd130, 8'd74, 8'd162, 8'd101, 8'd93, 8'd101, 8'd173, 8'd142, 8'd134, 8'd143, 8'd129, 8'd96, 8'd127, 8'd103, 8'd118, 8'd155, 8'd107, 8'd61, 8'd123, 8'd111, 8'd131, 8'd165, 8'd88, 8'd150, 8'd187, 8'd87, 8'd89, 8'd107, 8'd129, 8'd118, 8'd98, 8'd126, 8'd90, 8'd114, 8'd183, 8'd96, 8'd141, 8'd158, 8'd168, 8'd181, 8'd147, 8'd181, 8'd185, 8'd153, 8'd118, 8'd154, 8'd131, 8'd143, 8'd91, 8'd123, 8'd111, 8'd146, 8'd118, 8'd86, 8'd147, 8'd135, 8'd169, 8'd120, 8'd137, 8'd107, 8'd163, 8'd154, 8'd176, 8'd163, 8'd107, 8'd145, 8'd151, 8'd177, 8'd154, 8'd168, 8'd180, 8'd127, 8'd161, 8'd172, 8'd113, 8'd152, 8'd97, 8'd79, 8'd165, 8'd146, 8'd120, 8'd145, 8'd112, 8'd146, 8'd99, 8'd160, 8'd120, 8'd88, 8'd161, 8'd100, 8'd125, 8'd108, 8'd73, 8'd92, 8'd182, 8'd104, 8'd162, 8'd192, 8'd193, 8'd138, 8'd161, 8'd127, 8'd162, 8'd115, 8'd154, 8'd112, 8'd99, 8'd170, 8'd160, 8'd163, 8'd79, 8'd170, 8'd77, 8'd149, 8'd96, 8'd165, 8'd143, 8'd145, 8'd156, 8'd144, 8'd123, 8'd99, 8'd151, 8'd158, 8'd95, 8'd107, 8'd119, 8'd140, 8'd124, 8'd108, 8'd107, 8'd146, 8'd107, 8'd124, 8'd66, 8'd130, 8'd130, 8'd150, 8'd98, 8'd104, 8'd114, 8'd77, 8'd148, 8'd89, 8'd78, 8'd97, 8'd91, 8'd154, 8'd142, 8'd141, 8'd151, 8'd91, 8'd167, 8'd88, 8'd111, 8'd87, 8'd118, 8'd87, 8'd79, 8'd88, 8'd75, 8'd95, 8'd77, 8'd148, 8'd112, 8'd122, 8'd130, 8'd105, 8'd120, 8'd122, 8'd150, 8'd157, 8'd152})
) cell_0_74 (
    .clk(clk),
    .input_index(index_0_73_74),
    .input_value(value_0_73_74),
    .input_result(result_0_73_74),
    .input_enable(enable_0_73_74),
    .output_index(index_0_74_75),
    .output_value(value_0_74_75),
    .output_result(result_0_74_75),
    .output_enable(enable_0_74_75)
);

wire [10-1:0] index_0_75_76;
wire [`DATA_WIDTH-1:0] value_0_75_76;
wire [`DATA_WIDTH*4:0] result_0_75_76;
wire enable_0_75_76;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd103, 8'd82, 8'd165, 8'd116, 8'd95, 8'd95, 8'd133, 8'd145, 8'd89, 8'd60, 8'd119, 8'd49, 8'd144, 8'd107, 8'd102, 8'd84, 8'd81, 8'd132, 8'd132, 8'd78, 8'd152, 8'd69, 8'd149, 8'd152, 8'd76, 8'd83, 8'd108, 8'd95, 8'd137, 8'd146, 8'd73, 8'd103, 8'd104, 8'd108, 8'd103, 8'd130, 8'd125, 8'd70, 8'd75, 8'd154, 8'd125, 8'd95, 8'd159, 8'd92, 8'd88, 8'd74, 8'd135, 8'd164, 8'd159, 8'd149, 8'd165, 8'd112, 8'd107, 8'd136, 8'd153, 8'd143, 8'd161, 8'd94, 8'd161, 8'd175, 8'd184, 8'd157, 8'd122, 8'd174, 8'd172, 8'd99, 8'd86, 8'd151, 8'd119, 8'd111, 8'd76, 8'd59, 8'd96, 8'd54, 8'd87, 8'd96, 8'd53, 8'd75, 8'd89, 8'd108, 8'd59, 8'd95, 8'd84, 8'd156, 8'd131, 8'd92, 8'd116, 8'd132, 8'd119, 8'd165, 8'd119, 8'd132, 8'd148, 8'd98, 8'd109, 8'd65, 8'd156, 8'd60, 8'd76, 8'd82, 8'd138, 8'd120, 8'd134, 8'd97, 8'd117, 8'd123, 8'd43, 8'd48, 8'd65, 8'd122, 8'd99, 8'd143, 8'd111, 8'd79, 8'd162, 8'd167, 8'd82, 8'd165, 8'd142, 8'd135, 8'd121, 8'd79, 8'd81, 8'd156, 8'd95, 8'd121, 8'd75, 8'd69, 8'd76, 8'd145, 8'd92, 8'd73, 8'd77, 8'd90, 8'd60, 8'd111, 8'd89, 8'd90, 8'd81, 8'd124, 8'd128, 8'd147, 8'd120, 8'd94, 8'd78, 8'd89, 8'd107, 8'd114, 8'd159, 8'd93, 8'd166, 8'd94, 8'd119, 8'd154, 8'd127, 8'd66, 8'd153, 8'd61, 8'd103, 8'd143, 8'd107, 8'd102, 8'd87, 8'd162, 8'd109, 8'd126, 8'd103, 8'd107, 8'd137, 8'd107, 8'd154, 8'd148, 8'd107, 8'd117, 8'd136, 8'd79, 8'd112, 8'd127, 8'd113, 8'd131, 8'd112, 8'd152, 8'd129, 8'd140, 8'd108, 8'd161, 8'd157, 8'd144, 8'd93, 8'd155, 8'd110, 8'd133, 8'd99, 8'd117, 8'd165, 8'd148, 8'd127, 8'd134, 8'd104, 8'd107, 8'd78, 8'd125, 8'd105, 8'd118, 8'd158, 8'd161, 8'd105, 8'd83, 8'd106, 8'd154, 8'd114, 8'd118, 8'd113, 8'd112, 8'd154, 8'd146, 8'd89, 8'd112, 8'd136, 8'd92, 8'd109, 8'd106, 8'd126, 8'd102, 8'd80, 8'd47, 8'd123, 8'd62, 8'd161, 8'd116, 8'd121, 8'd145, 8'd96, 8'd95, 8'd144, 8'd66, 8'd162, 8'd82, 8'd110, 8'd170, 8'd102, 8'd172, 8'd128, 8'd146, 8'd81, 8'd113, 8'd74, 8'd46, 8'd64, 8'd118, 8'd119, 8'd115, 8'd128, 8'd60, 8'd63, 8'd117, 8'd112, 8'd83, 8'd151, 8'd149, 8'd138, 8'd64, 8'd53, 8'd57, 8'd116, 8'd183, 8'd168, 8'd155, 8'd144, 8'd91, 8'd104, 8'd160, 8'd164, 8'd96, 8'd126, 8'd67, 8'd125, 8'd105, 8'd130, 8'd108, 8'd80, 8'd40, 8'd45, 8'd104, 8'd129, 8'd112, 8'd96, 8'd59, 8'd78, 8'd145, 8'd46, 8'd114, 8'd129, 8'd112, 8'd158, 8'd96, 8'd112, 8'd128, 8'd136, 8'd134, 8'd128, 8'd60, 8'd73, 8'd88, 8'd103, 8'd125, 8'd81, 8'd96, 8'd141, 8'd35, 8'd76, 8'd115, 8'd143, 8'd131, 8'd61, 8'd127, 8'd130, 8'd91, 8'd134, 8'd155, 8'd148, 8'd183, 8'd147, 8'd161, 8'd164, 8'd79, 8'd68, 8'd133, 8'd135, 8'd79, 8'd37, 8'd87, 8'd137, 8'd81, 8'd100, 8'd124, 8'd112, 8'd103, 8'd104, 8'd137, 8'd133, 8'd136, 8'd63, 8'd61, 8'd69, 8'd69, 8'd133, 8'd142, 8'd101, 8'd198, 8'd170, 8'd184, 8'd138, 8'd132, 8'd157, 8'd96, 8'd112, 8'd143, 8'd66, 8'd56, 8'd71, 8'd82, 8'd88, 8'd121, 8'd139, 8'd119, 8'd103, 8'd126, 8'd103, 8'd94, 8'd131, 8'd94, 8'd127, 8'd57, 8'd89, 8'd175, 8'd176, 8'd167, 8'd181, 8'd187, 8'd93, 8'd87, 8'd65, 8'd140, 8'd97, 8'd168, 8'd98, 8'd134, 8'd88, 8'd121, 8'd159, 8'd78, 8'd135, 8'd49, 8'd130, 8'd59, 8'd145, 8'd80, 8'd90, 8'd157, 8'd132, 8'd97, 8'd134, 8'd98, 8'd183, 8'd118, 8'd148, 8'd160, 8'd130, 8'd153, 8'd129, 8'd122, 8'd176, 8'd152, 8'd145, 8'd103, 8'd144, 8'd130, 8'd118, 8'd83, 8'd72, 8'd98, 8'd100, 8'd143, 8'd104, 8'd150, 8'd111, 8'd100, 8'd64, 8'd86, 8'd87, 8'd69, 8'd106, 8'd117, 8'd223, 8'd124, 8'd113, 8'd149, 8'd118, 8'd109, 8'd135, 8'd120, 8'd146, 8'd149, 8'd72, 8'd90, 8'd91, 8'd82, 8'd141, 8'd126, 8'd184, 8'd190, 8'd116, 8'd100, 8'd101, 8'd58, 8'd19, 8'd81, 8'd80, 8'd125, 8'd129, 8'd196, 8'd175, 8'd166, 8'd152, 8'd197, 8'd113, 8'd176, 8'd207, 8'd194, 8'd122, 8'd96, 8'd116, 8'd70, 8'd57, 8'd103, 8'd163, 8'd187, 8'd235, 8'd222, 8'd141, 8'd161, 8'd129, 8'd66, 8'd83, 8'd74, 8'd74, 8'd122, 8'd101, 8'd120, 8'd169, 8'd212, 8'd211, 8'd173, 8'd174, 8'd169, 8'd184, 8'd100, 8'd77, 8'd50, 8'd46, 8'd48, 8'd155, 8'd160, 8'd85, 8'd190, 8'd166, 8'd156, 8'd148, 8'd102, 8'd116, 8'd48, 8'd79, 8'd33, 8'd63, 8'd36, 8'd22, 8'd105, 8'd148, 8'd186, 8'd99, 8'd176, 8'd138, 8'd135, 8'd116, 8'd92, 8'd72, 8'd52, 8'd80, 8'd129, 8'd62, 8'd80, 8'd110, 8'd115, 8'd222, 8'd222, 8'd200, 8'd166, 8'd91, 8'd70, 8'd80, 8'd69, 8'd79, 8'd80, 8'd63, 8'd60, 8'd67, 8'd120, 8'd132, 8'd143, 8'd68, 8'd138, 8'd125, 8'd123, 8'd129, 8'd53, 8'd129, 8'd139, 8'd59, 8'd139, 8'd118, 8'd195, 8'd153, 8'd140, 8'd183, 8'd154, 8'd149, 8'd130, 8'd97, 8'd134, 8'd61, 8'd103, 8'd109, 8'd100, 8'd51, 8'd71, 8'd65, 8'd143, 8'd86, 8'd119, 8'd71, 8'd93, 8'd55, 8'd99, 8'd103, 8'd93, 8'd86, 8'd91, 8'd85, 8'd169, 8'd164, 8'd224, 8'd199, 8'd165, 8'd127, 8'd144, 8'd159, 8'd106, 8'd86, 8'd63, 8'd58, 8'd109, 8'd87, 8'd146, 8'd82, 8'd110, 8'd72, 8'd55, 8'd62, 8'd71, 8'd107, 8'd53, 8'd45, 8'd153, 8'd66, 8'd129, 8'd153, 8'd116, 8'd188, 8'd152, 8'd161, 8'd141, 8'd125, 8'd129, 8'd152, 8'd105, 8'd165, 8'd149, 8'd131, 8'd83, 8'd151, 8'd121, 8'd106, 8'd121, 8'd73, 8'd141, 8'd106, 8'd84, 8'd60, 8'd78, 8'd107, 8'd73, 8'd89, 8'd85, 8'd98, 8'd129, 8'd144, 8'd113, 8'd133, 8'd200, 8'd178, 8'd179, 8'd148, 8'd116, 8'd150, 8'd119, 8'd118, 8'd112, 8'd116, 8'd146, 8'd57, 8'd67, 8'd60, 8'd110, 8'd134, 8'd102, 8'd56, 8'd84, 8'd103, 8'd95, 8'd120, 8'd129, 8'd79, 8'd135, 8'd122, 8'd86, 8'd172, 8'd194, 8'd122, 8'd161, 8'd133, 8'd114, 8'd123, 8'd149, 8'd86, 8'd135, 8'd67, 8'd133, 8'd118, 8'd141, 8'd134, 8'd123, 8'd163, 8'd111, 8'd110, 8'd126, 8'd103, 8'd105, 8'd141, 8'd120, 8'd132, 8'd103, 8'd100, 8'd93, 8'd148, 8'd98, 8'd187, 8'd170, 8'd163, 8'd124, 8'd142, 8'd79, 8'd145, 8'd140, 8'd106, 8'd88, 8'd114, 8'd149, 8'd167, 8'd157, 8'd92, 8'd164, 8'd126, 8'd113, 8'd85, 8'd99, 8'd102, 8'd88, 8'd155, 8'd149, 8'd91, 8'd159, 8'd126, 8'd93, 8'd142, 8'd125, 8'd93, 8'd143, 8'd103, 8'd58, 8'd147, 8'd136, 8'd129, 8'd155, 8'd85, 8'd125, 8'd115, 8'd86, 8'd113, 8'd133, 8'd86, 8'd167, 8'd137, 8'd130, 8'd158, 8'd143, 8'd132, 8'd110, 8'd79, 8'd95, 8'd92, 8'd91, 8'd145, 8'd101, 8'd166, 8'd150, 8'd118, 8'd95, 8'd112, 8'd125, 8'd77, 8'd103, 8'd95, 8'd151, 8'd166, 8'd100, 8'd114, 8'd109, 8'd83, 8'd128, 8'd104, 8'd94, 8'd101, 8'd133})
) cell_0_75 (
    .clk(clk),
    .input_index(index_0_74_75),
    .input_value(value_0_74_75),
    .input_result(result_0_74_75),
    .input_enable(enable_0_74_75),
    .output_index(index_0_75_76),
    .output_value(value_0_75_76),
    .output_result(result_0_75_76),
    .output_enable(enable_0_75_76)
);

wire [10-1:0] index_0_76_77;
wire [`DATA_WIDTH-1:0] value_0_76_77;
wire [`DATA_WIDTH*4:0] result_0_76_77;
wire enable_0_76_77;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd111, 8'd100, 8'd105, 8'd88, 8'd152, 8'd134, 8'd129, 8'd132, 8'd136, 8'd118, 8'd152, 8'd189, 8'd118, 8'd176, 8'd147, 8'd147, 8'd152, 8'd105, 8'd157, 8'd155, 8'd149, 8'd164, 8'd162, 8'd153, 8'd101, 8'd110, 8'd134, 8'd109, 8'd98, 8'd91, 8'd78, 8'd117, 8'd105, 8'd127, 8'd87, 8'd167, 8'd151, 8'd186, 8'd118, 8'd164, 8'd205, 8'd132, 8'd155, 8'd137, 8'd161, 8'd170, 8'd183, 8'd116, 8'd113, 8'd119, 8'd139, 8'd87, 8'd98, 8'd132, 8'd95, 8'd77, 8'd104, 8'd142, 8'd131, 8'd126, 8'd85, 8'd144, 8'd178, 8'd125, 8'd120, 8'd128, 8'd194, 8'd149, 8'd171, 8'd134, 8'd211, 8'd211, 8'd188, 8'd155, 8'd115, 8'd132, 8'd122, 8'd105, 8'd188, 8'd132, 8'd114, 8'd131, 8'd162, 8'd100, 8'd77, 8'd121, 8'd137, 8'd94, 8'd135, 8'd140, 8'd137, 8'd119, 8'd178, 8'd109, 8'd132, 8'd195, 8'd147, 8'd130, 8'd119, 8'd119, 8'd216, 8'd162, 8'd194, 8'd200, 8'd147, 8'd142, 8'd167, 8'd116, 8'd139, 8'd68, 8'd129, 8'd157, 8'd162, 8'd73, 8'd93, 8'd118, 8'd159, 8'd113, 8'd163, 8'd109, 8'd134, 8'd129, 8'd86, 8'd167, 8'd95, 8'd122, 8'd160, 8'd188, 8'd170, 8'd142, 8'd117, 8'd159, 8'd108, 8'd126, 8'd135, 8'd90, 8'd160, 8'd157, 8'd116, 8'd144, 8'd116, 8'd82, 8'd158, 8'd92, 8'd91, 8'd107, 8'd147, 8'd89, 8'd74, 8'd107, 8'd120, 8'd134, 8'd118, 8'd160, 8'd143, 8'd157, 8'd143, 8'd81, 8'd139, 8'd64, 8'd59, 8'd50, 8'd65, 8'd110, 8'd115, 8'd95, 8'd120, 8'd148, 8'd122, 8'd138, 8'd109, 8'd114, 8'd90, 8'd117, 8'd61, 8'd88, 8'd108, 8'd75, 8'd107, 8'd92, 8'd120, 8'd75, 8'd152, 8'd164, 8'd129, 8'd68, 8'd64, 8'd81, 8'd106, 8'd55, 8'd95, 8'd107, 8'd54, 8'd99, 8'd153, 8'd148, 8'd137, 8'd107, 8'd107, 8'd176, 8'd115, 8'd76, 8'd115, 8'd129, 8'd81, 8'd69, 8'd94, 8'd109, 8'd117, 8'd144, 8'd95, 8'd98, 8'd110, 8'd110, 8'd123, 8'd141, 8'd66, 8'd102, 8'd91, 8'd81, 8'd99, 8'd95, 8'd117, 8'd117, 8'd111, 8'd97, 8'd120, 8'd149, 8'd95, 8'd89, 8'd146, 8'd131, 8'd115, 8'd153, 8'd116, 8'd90, 8'd112, 8'd108, 8'd76, 8'd130, 8'd124, 8'd111, 8'd111, 8'd112, 8'd102, 8'd131, 8'd103, 8'd149, 8'd56, 8'd88, 8'd95, 8'd91, 8'd120, 8'd143, 8'd98, 8'd122, 8'd149, 8'd147, 8'd141, 8'd92, 8'd126, 8'd127, 8'd125, 8'd175, 8'd163, 8'd110, 8'd72, 8'd111, 8'd129, 8'd120, 8'd62, 8'd147, 8'd109, 8'd108, 8'd158, 8'd129, 8'd82, 8'd123, 8'd100, 8'd136, 8'd100, 8'd96, 8'd160, 8'd144, 8'd86, 8'd88, 8'd73, 8'd118, 8'd99, 8'd153, 8'd174, 8'd194, 8'd131, 8'd152, 8'd141, 8'd147, 8'd141, 8'd104, 8'd63, 8'd140, 8'd157, 8'd153, 8'd110, 8'd75, 8'd119, 8'd140, 8'd154, 8'd129, 8'd169, 8'd154, 8'd69, 8'd98, 8'd122, 8'd108, 8'd103, 8'd142, 8'd136, 8'd156, 8'd169, 8'd170, 8'd154, 8'd94, 8'd94, 8'd82, 8'd103, 8'd124, 8'd94, 8'd76, 8'd119, 8'd142, 8'd88, 8'd155, 8'd67, 8'd64, 8'd68, 8'd160, 8'd99, 8'd98, 8'd72, 8'd133, 8'd111, 8'd130, 8'd163, 8'd196, 8'd168, 8'd224, 8'd209, 8'd113, 8'd139, 8'd98, 8'd89, 8'd115, 8'd158, 8'd164, 8'd130, 8'd76, 8'd105, 8'd117, 8'd95, 8'd86, 8'd113, 8'd147, 8'd103, 8'd94, 8'd108, 8'd110, 8'd82, 8'd101, 8'd87, 8'd139, 8'd119, 8'd150, 8'd145, 8'd198, 8'd199, 8'd203, 8'd140, 8'd60, 8'd83, 8'd69, 8'd109, 8'd161, 8'd76, 8'd154, 8'd159, 8'd115, 8'd142, 8'd183, 8'd163, 8'd150, 8'd109, 8'd168, 8'd132, 8'd168, 8'd94, 8'd96, 8'd86, 8'd75, 8'd156, 8'd166, 8'd173, 8'd165, 8'd130, 8'd129, 8'd155, 8'd124, 8'd126, 8'd161, 8'd105, 8'd108, 8'd149, 8'd86, 8'd114, 8'd96, 8'd182, 8'd135, 8'd137, 8'd141, 8'd83, 8'd73, 8'd145, 8'd125, 8'd167, 8'd66, 8'd92, 8'd138, 8'd127, 8'd144, 8'd129, 8'd137, 8'd153, 8'd171, 8'd148, 8'd96, 8'd127, 8'd156, 8'd164, 8'd151, 8'd168, 8'd116, 8'd146, 8'd132, 8'd115, 8'd196, 8'd130, 8'd124, 8'd95, 8'd89, 8'd124, 8'd137, 8'd112, 8'd119, 8'd152, 8'd91, 8'd136, 8'd167, 8'd186, 8'd186, 8'd198, 8'd101, 8'd86, 8'd69, 8'd60, 8'd137, 8'd147, 8'd171, 8'd154, 8'd175, 8'd102, 8'd189, 8'd117, 8'd165, 8'd148, 8'd167, 8'd126, 8'd108, 8'd169, 8'd200, 8'd189, 8'd150, 8'd92, 8'd113, 8'd148, 8'd107, 8'd138, 8'd193, 8'd160, 8'd161, 8'd127, 8'd66, 8'd109, 8'd134, 8'd183, 8'd164, 8'd156, 8'd186, 8'd196, 8'd180, 8'd176, 8'd97, 8'd153, 8'd124, 8'd138, 8'd96, 8'd79, 8'd107, 8'd175, 8'd203, 8'd133, 8'd146, 8'd155, 8'd116, 8'd142, 8'd183, 8'd173, 8'd161, 8'd109, 8'd157, 8'd142, 8'd162, 8'd122, 8'd124, 8'd127, 8'd159, 8'd147, 8'd193, 8'd151, 8'd163, 8'd171, 8'd138, 8'd135, 8'd113, 8'd102, 8'd132, 8'd126, 8'd130, 8'd131, 8'd118, 8'd182, 8'd158, 8'd178, 8'd133, 8'd174, 8'd172, 8'd131, 8'd86, 8'd177, 8'd128, 8'd195, 8'd176, 8'd139, 8'd200, 8'd147, 8'd119, 8'd160, 8'd104, 8'd92, 8'd129, 8'd103, 8'd69, 8'd146, 8'd107, 8'd188, 8'd186, 8'd139, 8'd98, 8'd91, 8'd134, 8'd175, 8'd105, 8'd114, 8'd190, 8'd97, 8'd142, 8'd176, 8'd171, 8'd164, 8'd193, 8'd166, 8'd214, 8'd127, 8'd137, 8'd147, 8'd108, 8'd131, 8'd127, 8'd98, 8'd131, 8'd152, 8'd132, 8'd174, 8'd174, 8'd98, 8'd99, 8'd127, 8'd149, 8'd77, 8'd155, 8'd163, 8'd95, 8'd157, 8'd93, 8'd105, 8'd150, 8'd158, 8'd116, 8'd148, 8'd183, 8'd144, 8'd97, 8'd90, 8'd108, 8'd116, 8'd107, 8'd164, 8'd154, 8'd147, 8'd110, 8'd155, 8'd113, 8'd68, 8'd137, 8'd59, 8'd131, 8'd142, 8'd92, 8'd127, 8'd79, 8'd71, 8'd154, 8'd99, 8'd106, 8'd139, 8'd159, 8'd119, 8'd99, 8'd117, 8'd104, 8'd77, 8'd114, 8'd145, 8'd71, 8'd81, 8'd108, 8'd149, 8'd75, 8'd163, 8'd106, 8'd155, 8'd114, 8'd85, 8'd131, 8'd79, 8'd125, 8'd139, 8'd103, 8'd119, 8'd56, 8'd53, 8'd92, 8'd128, 8'd76, 8'd126, 8'd58, 8'd107, 8'd141, 8'd105, 8'd114, 8'd108, 8'd112, 8'd157, 8'd93, 8'd117, 8'd106, 8'd168, 8'd75, 8'd118, 8'd120, 8'd104, 8'd160, 8'd117, 8'd162, 8'd134, 8'd85, 8'd121, 8'd77, 8'd137, 8'd60, 8'd65, 8'd90, 8'd92, 8'd145, 8'd108, 8'd102, 8'd91, 8'd85, 8'd102, 8'd160, 8'd95, 8'd88, 8'd135, 8'd113, 8'd148, 8'd145, 8'd93, 8'd138, 8'd88, 8'd100, 8'd126, 8'd111, 8'd96, 8'd55, 8'd121, 8'd52, 8'd42, 8'd57, 8'd119, 8'd59, 8'd137, 8'd105, 8'd126, 8'd115, 8'd131, 8'd126, 8'd70, 8'd70, 8'd124, 8'd85, 8'd104, 8'd135, 8'd147, 8'd129, 8'd117, 8'd111, 8'd93, 8'd123, 8'd97, 8'd52, 8'd73, 8'd102, 8'd114, 8'd70, 8'd125, 8'd105, 8'd110, 8'd82, 8'd120, 8'd71, 8'd70, 8'd113, 8'd155, 8'd105, 8'd135, 8'd118, 8'd153, 8'd156, 8'd111, 8'd78, 8'd90, 8'd80, 8'd137, 8'd94, 8'd121, 8'd165, 8'd157, 8'd78, 8'd163, 8'd153, 8'd69, 8'd143, 8'd68, 8'd145, 8'd143, 8'd73, 8'd109, 8'd75, 8'd118, 8'd155, 8'd96, 8'd87, 8'd166, 8'd78, 8'd121, 8'd162})
) cell_0_76 (
    .clk(clk),
    .input_index(index_0_75_76),
    .input_value(value_0_75_76),
    .input_result(result_0_75_76),
    .input_enable(enable_0_75_76),
    .output_index(index_0_76_77),
    .output_value(value_0_76_77),
    .output_result(result_0_76_77),
    .output_enable(enable_0_76_77)
);

wire [10-1:0] index_0_77_78;
wire [`DATA_WIDTH-1:0] value_0_77_78;
wire [`DATA_WIDTH*4:0] result_0_77_78;
wire enable_0_77_78;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd135, 8'd148, 8'd76, 8'd83, 8'd72, 8'd84, 8'd146, 8'd97, 8'd114, 8'd80, 8'd125, 8'd152, 8'd57, 8'd135, 8'd126, 8'd140, 8'd121, 8'd64, 8'd80, 8'd67, 8'd132, 8'd112, 8'd134, 8'd162, 8'd136, 8'd103, 8'd118, 8'd86, 8'd142, 8'd167, 8'd124, 8'd145, 8'd142, 8'd103, 8'd83, 8'd129, 8'd109, 8'd137, 8'd86, 8'd56, 8'd66, 8'd119, 8'd69, 8'd84, 8'd107, 8'd52, 8'd84, 8'd109, 8'd59, 8'd80, 8'd85, 8'd97, 8'd141, 8'd82, 8'd129, 8'd96, 8'd105, 8'd93, 8'd154, 8'd101, 8'd97, 8'd138, 8'd62, 8'd124, 8'd151, 8'd154, 8'd93, 8'd84, 8'd84, 8'd77, 8'd148, 8'd168, 8'd161, 8'd116, 8'd119, 8'd87, 8'd110, 8'd159, 8'd153, 8'd122, 8'd127, 8'd83, 8'd85, 8'd80, 8'd86, 8'd80, 8'd176, 8'd115, 8'd124, 8'd158, 8'd69, 8'd133, 8'd131, 8'd150, 8'd172, 8'd178, 8'd106, 8'd146, 8'd152, 8'd182, 8'd170, 8'd106, 8'd168, 8'd124, 8'd162, 8'd102, 8'd89, 8'd98, 8'd136, 8'd131, 8'd91, 8'd88, 8'd117, 8'd157, 8'd96, 8'd112, 8'd98, 8'd158, 8'd86, 8'd128, 8'd97, 8'd94, 8'd160, 8'd149, 8'd103, 8'd180, 8'd154, 8'd174, 8'd113, 8'd155, 8'd141, 8'd126, 8'd100, 8'd138, 8'd156, 8'd165, 8'd141, 8'd150, 8'd80, 8'd164, 8'd78, 8'd118, 8'd133, 8'd119, 8'd110, 8'd121, 8'd126, 8'd135, 8'd116, 8'd113, 8'd115, 8'd142, 8'd115, 8'd84, 8'd117, 8'd96, 8'd95, 8'd126, 8'd104, 8'd87, 8'd97, 8'd87, 8'd175, 8'd151, 8'd179, 8'd118, 8'd135, 8'd74, 8'd162, 8'd149, 8'd145, 8'd105, 8'd150, 8'd156, 8'd139, 8'd156, 8'd169, 8'd126, 8'd143, 8'd161, 8'd177, 8'd148, 8'd95, 8'd103, 8'd106, 8'd95, 8'd162, 8'd103, 8'd140, 8'd170, 8'd161, 8'd169, 8'd130, 8'd180, 8'd127, 8'd139, 8'd97, 8'd122, 8'd168, 8'd92, 8'd158, 8'd149, 8'd118, 8'd126, 8'd100, 8'd180, 8'd102, 8'd141, 8'd157, 8'd106, 8'd94, 8'd98, 8'd82, 8'd141, 8'd146, 8'd122, 8'd112, 8'd201, 8'd128, 8'd179, 8'd194, 8'd144, 8'd104, 8'd105, 8'd84, 8'd101, 8'd121, 8'd152, 8'd173, 8'd185, 8'd106, 8'd98, 8'd97, 8'd96, 8'd159, 8'd105, 8'd125, 8'd89, 8'd73, 8'd128, 8'd153, 8'd97, 8'd149, 8'd144, 8'd134, 8'd166, 8'd206, 8'd191, 8'd199, 8'd152, 8'd131, 8'd90, 8'd153, 8'd139, 8'd96, 8'd103, 8'd133, 8'd123, 8'd197, 8'd139, 8'd95, 8'd145, 8'd169, 8'd100, 8'd104, 8'd68, 8'd89, 8'd74, 8'd71, 8'd155, 8'd104, 8'd111, 8'd170, 8'd175, 8'd117, 8'd174, 8'd139, 8'd122, 8'd162, 8'd121, 8'd138, 8'd160, 8'd184, 8'd182, 8'd167, 8'd181, 8'd160, 8'd84, 8'd181, 8'd160, 8'd104, 8'd127, 8'd72, 8'd128, 8'd103, 8'd56, 8'd78, 8'd69, 8'd139, 8'd80, 8'd126, 8'd181, 8'd170, 8'd139, 8'd158, 8'd120, 8'd134, 8'd109, 8'd107, 8'd153, 8'd128, 8'd119, 8'd139, 8'd152, 8'd132, 8'd133, 8'd109, 8'd86, 8'd112, 8'd79, 8'd61, 8'd96, 8'd80, 8'd152, 8'd80, 8'd67, 8'd114, 8'd95, 8'd96, 8'd80, 8'd98, 8'd163, 8'd104, 8'd94, 8'd176, 8'd88, 8'd154, 8'd119, 8'd166, 8'd166, 8'd146, 8'd100, 8'd102, 8'd145, 8'd147, 8'd147, 8'd120, 8'd133, 8'd103, 8'd119, 8'd152, 8'd102, 8'd102, 8'd126, 8'd101, 8'd88, 8'd138, 8'd116, 8'd141, 8'd159, 8'd147, 8'd157, 8'd139, 8'd128, 8'd123, 8'd122, 8'd164, 8'd139, 8'd154, 8'd77, 8'd119, 8'd133, 8'd67, 8'd79, 8'd118, 8'd75, 8'd77, 8'd164, 8'd169, 8'd172, 8'd129, 8'd136, 8'd131, 8'd79, 8'd82, 8'd50, 8'd73, 8'd95, 8'd71, 8'd147, 8'd165, 8'd161, 8'd143, 8'd136, 8'd102, 8'd106, 8'd61, 8'd62, 8'd88, 8'd110, 8'd148, 8'd95, 8'd119, 8'd96, 8'd70, 8'd161, 8'd179, 8'd152, 8'd139, 8'd82, 8'd147, 8'd87, 8'd74, 8'd48, 8'd66, 8'd90, 8'd101, 8'd139, 8'd130, 8'd76, 8'd126, 8'd113, 8'd138, 8'd71, 8'd138, 8'd82, 8'd43, 8'd86, 8'd125, 8'd83, 8'd93, 8'd119, 8'd77, 8'd173, 8'd100, 8'd165, 8'd146, 8'd90, 8'd58, 8'd108, 8'd110, 8'd81, 8'd107, 8'd83, 8'd114, 8'd90, 8'd101, 8'd128, 8'd77, 8'd182, 8'd149, 8'd136, 8'd138, 8'd80, 8'd125, 8'd168, 8'd148, 8'd156, 8'd87, 8'd67, 8'd133, 8'd162, 8'd158, 8'd140, 8'd81, 8'd113, 8'd128, 8'd48, 8'd85, 8'd104, 8'd68, 8'd111, 8'd137, 8'd154, 8'd124, 8'd114, 8'd178, 8'd115, 8'd180, 8'd202, 8'd118, 8'd99, 8'd178, 8'd135, 8'd129, 8'd129, 8'd148, 8'd97, 8'd137, 8'd80, 8'd90, 8'd108, 8'd62, 8'd98, 8'd116, 8'd126, 8'd95, 8'd94, 8'd122, 8'd138, 8'd188, 8'd137, 8'd102, 8'd102, 8'd111, 8'd202, 8'd158, 8'd141, 8'd166, 8'd178, 8'd149, 8'd143, 8'd93, 8'd143, 8'd161, 8'd165, 8'd105, 8'd150, 8'd130, 8'd147, 8'd70, 8'd105, 8'd65, 8'd142, 8'd140, 8'd143, 8'd98, 8'd175, 8'd83, 8'd80, 8'd92, 8'd66, 8'd174, 8'd160, 8'd152, 8'd169, 8'd119, 8'd113, 8'd161, 8'd120, 8'd127, 8'd167, 8'd149, 8'd140, 8'd113, 8'd89, 8'd87, 8'd136, 8'd164, 8'd89, 8'd148, 8'd106, 8'd159, 8'd96, 8'd110, 8'd183, 8'd138, 8'd145, 8'd80, 8'd143, 8'd85, 8'd173, 8'd190, 8'd138, 8'd163, 8'd86, 8'd140, 8'd171, 8'd105, 8'd118, 8'd90, 8'd97, 8'd170, 8'd177, 8'd94, 8'd132, 8'd99, 8'd146, 8'd146, 8'd94, 8'd184, 8'd97, 8'd187, 8'd178, 8'd106, 8'd135, 8'd94, 8'd143, 8'd168, 8'd106, 8'd110, 8'd135, 8'd69, 8'd136, 8'd148, 8'd145, 8'd130, 8'd90, 8'd87, 8'd115, 8'd85, 8'd170, 8'd140, 8'd133, 8'd102, 8'd137, 8'd141, 8'd102, 8'd171, 8'd143, 8'd144, 8'd94, 8'd99, 8'd153, 8'd122, 8'd96, 8'd142, 8'd153, 8'd98, 8'd60, 8'd92, 8'd68, 8'd140, 8'd111, 8'd88, 8'd124, 8'd104, 8'd110, 8'd97, 8'd138, 8'd101, 8'd78, 8'd144, 8'd140, 8'd144, 8'd115, 8'd91, 8'd114, 8'd148, 8'd86, 8'd165, 8'd126, 8'd150, 8'd162, 8'd164, 8'd146, 8'd143, 8'd139, 8'd92, 8'd112, 8'd89, 8'd77, 8'd119, 8'd161, 8'd100, 8'd110, 8'd161, 8'd117, 8'd181, 8'd162, 8'd168, 8'd122, 8'd109, 8'd169, 8'd141, 8'd117, 8'd159, 8'd84, 8'd117, 8'd171, 8'd131, 8'd129, 8'd124, 8'd71, 8'd151, 8'd136, 8'd92, 8'd73, 8'd54, 8'd87, 8'd64, 8'd94, 8'd170, 8'd143, 8'd126, 8'd172, 8'd169, 8'd153, 8'd141, 8'd102, 8'd155, 8'd173, 8'd138, 8'd74, 8'd117, 8'd78, 8'd148, 8'd105, 8'd145, 8'd114, 8'd151, 8'd131, 8'd162, 8'd88, 8'd58, 8'd96, 8'd123, 8'd57, 8'd80, 8'd79, 8'd66, 8'd166, 8'd131, 8'd116, 8'd96, 8'd105, 8'd136, 8'd99, 8'd63, 8'd147, 8'd89, 8'd96, 8'd116, 8'd144, 8'd109, 8'd110, 8'd97, 8'd128, 8'd154, 8'd128, 8'd166, 8'd154, 8'd179, 8'd104, 8'd94, 8'd102, 8'd70, 8'd88, 8'd133, 8'd102, 8'd87, 8'd100, 8'd133, 8'd114, 8'd156, 8'd93, 8'd85, 8'd123, 8'd155, 8'd78, 8'd112, 8'd115, 8'd138, 8'd90, 8'd116, 8'd93, 8'd78, 8'd73, 8'd99, 8'd158, 8'd105, 8'd129, 8'd75, 8'd122, 8'd130, 8'd118, 8'd87, 8'd160, 8'd161, 8'd89, 8'd156, 8'd139, 8'd90, 8'd160, 8'd139, 8'd114, 8'd112, 8'd98, 8'd82, 8'd144, 8'd117, 8'd108, 8'd110, 8'd114})
) cell_0_77 (
    .clk(clk),
    .input_index(index_0_76_77),
    .input_value(value_0_76_77),
    .input_result(result_0_76_77),
    .input_enable(enable_0_76_77),
    .output_index(index_0_77_78),
    .output_value(value_0_77_78),
    .output_result(result_0_77_78),
    .output_enable(enable_0_77_78)
);

wire [10-1:0] index_0_78_79;
wire [`DATA_WIDTH-1:0] value_0_78_79;
wire [`DATA_WIDTH*4:0] result_0_78_79;
wire enable_0_78_79;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd83, 8'd96, 8'd112, 8'd137, 8'd123, 8'd116, 8'd69, 8'd116, 8'd113, 8'd81, 8'd64, 8'd123, 8'd112, 8'd160, 8'd46, 8'd66, 8'd93, 8'd112, 8'd122, 8'd146, 8'd88, 8'd118, 8'd86, 8'd158, 8'd71, 8'd80, 8'd146, 8'd72, 8'd117, 8'd88, 8'd101, 8'd165, 8'd72, 8'd152, 8'd162, 8'd106, 8'd148, 8'd155, 8'd149, 8'd131, 8'd174, 8'd164, 8'd80, 8'd87, 8'd124, 8'd115, 8'd121, 8'd125, 8'd124, 8'd80, 8'd97, 8'd110, 8'd135, 8'd85, 8'd103, 8'd163, 8'd160, 8'd150, 8'd85, 8'd85, 8'd77, 8'd100, 8'd132, 8'd174, 8'd92, 8'd97, 8'd173, 8'd154, 8'd148, 8'd77, 8'd63, 8'd70, 8'd145, 8'd133, 8'd95, 8'd61, 8'd53, 8'd104, 8'd103, 8'd109, 8'd86, 8'd76, 8'd79, 8'd111, 8'd88, 8'd78, 8'd104, 8'd107, 8'd128, 8'd136, 8'd149, 8'd104, 8'd97, 8'd122, 8'd73, 8'd122, 8'd149, 8'd142, 8'd88, 8'd78, 8'd138, 8'd96, 8'd92, 8'd95, 8'd61, 8'd121, 8'd49, 8'd35, 8'd90, 8'd163, 8'd95, 8'd140, 8'd145, 8'd100, 8'd74, 8'd149, 8'd177, 8'd163, 8'd105, 8'd148, 8'd120, 8'd136, 8'd137, 8'd131, 8'd97, 8'd95, 8'd163, 8'd122, 8'd114, 8'd92, 8'd134, 8'd160, 8'd105, 8'd108, 8'd114, 8'd119, 8'd151, 8'd82, 8'd130, 8'd156, 8'd79, 8'd70, 8'd80, 8'd92, 8'd159, 8'd93, 8'd168, 8'd144, 8'd107, 8'd135, 8'd99, 8'd140, 8'd137, 8'd154, 8'd177, 8'd142, 8'd97, 8'd136, 8'd148, 8'd118, 8'd169, 8'd127, 8'd108, 8'd109, 8'd87, 8'd136, 8'd71, 8'd128, 8'd111, 8'd154, 8'd99, 8'd154, 8'd164, 8'd149, 8'd110, 8'd134, 8'd165, 8'd192, 8'd178, 8'd141, 8'd85, 8'd101, 8'd193, 8'd138, 8'd183, 8'd130, 8'd86, 8'd112, 8'd119, 8'd154, 8'd92, 8'd116, 8'd124, 8'd117, 8'd134, 8'd90, 8'd136, 8'd156, 8'd140, 8'd164, 8'd145, 8'd183, 8'd98, 8'd188, 8'd183, 8'd119, 8'd153, 8'd117, 8'd115, 8'd151, 8'd109, 8'd199, 8'd132, 8'd148, 8'd129, 8'd125, 8'd190, 8'd95, 8'd114, 8'd80, 8'd99, 8'd101, 8'd68, 8'd170, 8'd166, 8'd150, 8'd213, 8'd147, 8'd166, 8'd204, 8'd160, 8'd139, 8'd158, 8'd184, 8'd122, 8'd122, 8'd166, 8'd98, 8'd116, 8'd115, 8'd216, 8'd118, 8'd196, 8'd117, 8'd100, 8'd104, 8'd67, 8'd141, 8'd57, 8'd123, 8'd62, 8'd92, 8'd97, 8'd148, 8'd177, 8'd169, 8'd148, 8'd173, 8'd190, 8'd164, 8'd150, 8'd158, 8'd183, 8'd96, 8'd114, 8'd167, 8'd122, 8'd120, 8'd215, 8'd207, 8'd121, 8'd109, 8'd121, 8'd141, 8'd159, 8'd158, 8'd111, 8'd150, 8'd105, 8'd96, 8'd172, 8'd109, 8'd204, 8'd120, 8'd98, 8'd151, 8'd84, 8'd179, 8'd136, 8'd84, 8'd158, 8'd156, 8'd87, 8'd92, 8'd182, 8'd192, 8'd213, 8'd140, 8'd182, 8'd161, 8'd159, 8'd153, 8'd117, 8'd119, 8'd119, 8'd78, 8'd73, 8'd84, 8'd87, 8'd108, 8'd139, 8'd134, 8'd96, 8'd93, 8'd141, 8'd63, 8'd77, 8'd103, 8'd127, 8'd119, 8'd155, 8'd109, 8'd186, 8'd115, 8'd163, 8'd191, 8'd101, 8'd157, 8'd94, 8'd171, 8'd131, 8'd153, 8'd119, 8'd126, 8'd149, 8'd86, 8'd149, 8'd123, 8'd174, 8'd174, 8'd91, 8'd115, 8'd122, 8'd118, 8'd136, 8'd109, 8'd140, 8'd87, 8'd116, 8'd109, 8'd148, 8'd184, 8'd104, 8'd100, 8'd130, 8'd138, 8'd78, 8'd110, 8'd89, 8'd82, 8'd150, 8'd58, 8'd141, 8'd74, 8'd155, 8'd160, 8'd142, 8'd166, 8'd124, 8'd81, 8'd107, 8'd151, 8'd122, 8'd70, 8'd161, 8'd162, 8'd113, 8'd190, 8'd177, 8'd111, 8'd150, 8'd93, 8'd62, 8'd57, 8'd134, 8'd100, 8'd131, 8'd98, 8'd152, 8'd79, 8'd77, 8'd99, 8'd107, 8'd106, 8'd197, 8'd148, 8'd150, 8'd137, 8'd108, 8'd148, 8'd139, 8'd151, 8'd152, 8'd111, 8'd91, 8'd101, 8'd127, 8'd138, 8'd100, 8'd69, 8'd50, 8'd128, 8'd92, 8'd96, 8'd72, 8'd88, 8'd87, 8'd81, 8'd130, 8'd120, 8'd166, 8'd92, 8'd190, 8'd225, 8'd148, 8'd161, 8'd161, 8'd149, 8'd105, 8'd93, 8'd140, 8'd111, 8'd129, 8'd118, 8'd101, 8'd102, 8'd137, 8'd126, 8'd53, 8'd130, 8'd65, 8'd54, 8'd56, 8'd114, 8'd132, 8'd71, 8'd132, 8'd82, 8'd128, 8'd78, 8'd101, 8'd138, 8'd116, 8'd144, 8'd178, 8'd124, 8'd70, 8'd52, 8'd96, 8'd100, 8'd112, 8'd66, 8'd80, 8'd80, 8'd50, 8'd66, 8'd130, 8'd157, 8'd118, 8'd138, 8'd90, 8'd147, 8'd90, 8'd80, 8'd111, 8'd73, 8'd99, 8'd119, 8'd119, 8'd62, 8'd117, 8'd80, 8'd99, 8'd69, 8'd70, 8'd114, 8'd55, 8'd104, 8'd57, 8'd140, 8'd86, 8'd148, 8'd104, 8'd94, 8'd103, 8'd159, 8'd172, 8'd83, 8'd81, 8'd139, 8'd89, 8'd88, 8'd96, 8'd71, 8'd118, 8'd119, 8'd108, 8'd96, 8'd140, 8'd118, 8'd105, 8'd77, 8'd65, 8'd89, 8'd68, 8'd122, 8'd163, 8'd117, 8'd136, 8'd111, 8'd160, 8'd93, 8'd157, 8'd97, 8'd171, 8'd84, 8'd95, 8'd109, 8'd154, 8'd54, 8'd137, 8'd78, 8'd146, 8'd70, 8'd137, 8'd137, 8'd136, 8'd54, 8'd104, 8'd103, 8'd113, 8'd75, 8'd110, 8'd98, 8'd136, 8'd136, 8'd155, 8'd161, 8'd155, 8'd133, 8'd139, 8'd143, 8'd166, 8'd172, 8'd148, 8'd107, 8'd86, 8'd91, 8'd94, 8'd131, 8'd125, 8'd124, 8'd97, 8'd142, 8'd79, 8'd68, 8'd72, 8'd96, 8'd118, 8'd61, 8'd141, 8'd164, 8'd125, 8'd119, 8'd109, 8'd156, 8'd128, 8'd161, 8'd168, 8'd89, 8'd151, 8'd156, 8'd158, 8'd162, 8'd127, 8'd149, 8'd138, 8'd116, 8'd122, 8'd159, 8'd118, 8'd100, 8'd49, 8'd116, 8'd104, 8'd62, 8'd121, 8'd123, 8'd88, 8'd98, 8'd127, 8'd110, 8'd136, 8'd163, 8'd100, 8'd158, 8'd88, 8'd107, 8'd78, 8'd159, 8'd101, 8'd129, 8'd122, 8'd71, 8'd84, 8'd72, 8'd166, 8'd113, 8'd118, 8'd124, 8'd64, 8'd56, 8'd149, 8'd93, 8'd148, 8'd162, 8'd169, 8'd113, 8'd169, 8'd186, 8'd144, 8'd183, 8'd109, 8'd105, 8'd180, 8'd92, 8'd133, 8'd87, 8'd157, 8'd140, 8'd101, 8'd79, 8'd81, 8'd93, 8'd98, 8'd92, 8'd130, 8'd89, 8'd101, 8'd115, 8'd90, 8'd104, 8'd146, 8'd153, 8'd172, 8'd118, 8'd179, 8'd170, 8'd133, 8'd101, 8'd171, 8'd164, 8'd195, 8'd150, 8'd157, 8'd174, 8'd110, 8'd84, 8'd141, 8'd131, 8'd68, 8'd136, 8'd89, 8'd147, 8'd162, 8'd159, 8'd165, 8'd188, 8'd153, 8'd112, 8'd132, 8'd156, 8'd193, 8'd168, 8'd199, 8'd152, 8'd212, 8'd215, 8'd177, 8'd137, 8'd152, 8'd161, 8'd113, 8'd179, 8'd173, 8'd93, 8'd129, 8'd163, 8'd165, 8'd125, 8'd92, 8'd99, 8'd166, 8'd151, 8'd160, 8'd163, 8'd133, 8'd137, 8'd144, 8'd132, 8'd201, 8'd193, 8'd154, 8'd226, 8'd223, 8'd215, 8'd171, 8'd133, 8'd151, 8'd176, 8'd170, 8'd134, 8'd162, 8'd142, 8'd164, 8'd141, 8'd103, 8'd168, 8'd112, 8'd164, 8'd82, 8'd103, 8'd81, 8'd109, 8'd117, 8'd141, 8'd140, 8'd109, 8'd186, 8'd183, 8'd119, 8'd159, 8'd166, 8'd126, 8'd158, 8'd169, 8'd185, 8'd122, 8'd161, 8'd154, 8'd128, 8'd153, 8'd93, 8'd77, 8'd80, 8'd143, 8'd163, 8'd100, 8'd147, 8'd147, 8'd123, 8'd163, 8'd152, 8'd120, 8'd80, 8'd155, 8'd167, 8'd75, 8'd93, 8'd98, 8'd166, 8'd110, 8'd129, 8'd163, 8'd78, 8'd92, 8'd170, 8'd165, 8'd118, 8'd148, 8'd110, 8'd138, 8'd80, 8'd105})
) cell_0_78 (
    .clk(clk),
    .input_index(index_0_77_78),
    .input_value(value_0_77_78),
    .input_result(result_0_77_78),
    .input_enable(enable_0_77_78),
    .output_index(index_0_78_79),
    .output_value(value_0_78_79),
    .output_result(result_0_78_79),
    .output_enable(enable_0_78_79)
);

wire [10-1:0] index_0_79_80;
wire [`DATA_WIDTH-1:0] value_0_79_80;
wire [`DATA_WIDTH*4:0] result_0_79_80;
wire enable_0_79_80;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd160, 8'd134, 8'd160, 8'd162, 8'd65, 8'd139, 8'd148, 8'd68, 8'd120, 8'd120, 8'd122, 8'd66, 8'd141, 8'd96, 8'd37, 8'd134, 8'd137, 8'd94, 8'd155, 8'd102, 8'd131, 8'd88, 8'd116, 8'd102, 8'd170, 8'd72, 8'd161, 8'd118, 8'd90, 8'd158, 8'd157, 8'd104, 8'd129, 8'd138, 8'd145, 8'd126, 8'd94, 8'd83, 8'd107, 8'd115, 8'd112, 8'd136, 8'd86, 8'd99, 8'd150, 8'd117, 8'd135, 8'd162, 8'd121, 8'd140, 8'd84, 8'd162, 8'd109, 8'd100, 8'd143, 8'd72, 8'd132, 8'd129, 8'd172, 8'd101, 8'd156, 8'd108, 8'd159, 8'd150, 8'd121, 8'd152, 8'd62, 8'd132, 8'd70, 8'd120, 8'd88, 8'd94, 8'd80, 8'd108, 8'd71, 8'd136, 8'd147, 8'd103, 8'd131, 8'd79, 8'd126, 8'd130, 8'd85, 8'd71, 8'd124, 8'd91, 8'd162, 8'd116, 8'd107, 8'd95, 8'd121, 8'd111, 8'd125, 8'd102, 8'd142, 8'd164, 8'd85, 8'd158, 8'd140, 8'd125, 8'd102, 8'd157, 8'd68, 8'd113, 8'd75, 8'd62, 8'd98, 8'd140, 8'd82, 8'd90, 8'd95, 8'd89, 8'd115, 8'd103, 8'd79, 8'd136, 8'd111, 8'd159, 8'd152, 8'd156, 8'd128, 8'd145, 8'd156, 8'd106, 8'd159, 8'd85, 8'd150, 8'd83, 8'd83, 8'd122, 8'd126, 8'd90, 8'd87, 8'd132, 8'd92, 8'd60, 8'd73, 8'd140, 8'd74, 8'd123, 8'd78, 8'd137, 8'd120, 8'd134, 8'd93, 8'd126, 8'd118, 8'd95, 8'd140, 8'd147, 8'd128, 8'd156, 8'd140, 8'd81, 8'd82, 8'd142, 8'd128, 8'd155, 8'd176, 8'd187, 8'd133, 8'd144, 8'd77, 8'd99, 8'd100, 8'd80, 8'd108, 8'd130, 8'd165, 8'd101, 8'd182, 8'd172, 8'd95, 8'd167, 8'd106, 8'd109, 8'd102, 8'd174, 8'd171, 8'd111, 8'd105, 8'd160, 8'd120, 8'd123, 8'd117, 8'd149, 8'd128, 8'd92, 8'd131, 8'd169, 8'd143, 8'd153, 8'd95, 8'd115, 8'd166, 8'd145, 8'd108, 8'd128, 8'd178, 8'd181, 8'd178, 8'd127, 8'd162, 8'd171, 8'd155, 8'd98, 8'd97, 8'd86, 8'd116, 8'd138, 8'd159, 8'd69, 8'd162, 8'd170, 8'd88, 8'd97, 8'd133, 8'd105, 8'd134, 8'd140, 8'd162, 8'd81, 8'd126, 8'd94, 8'd118, 8'd136, 8'd109, 8'd131, 8'd149, 8'd107, 8'd139, 8'd149, 8'd132, 8'd155, 8'd97, 8'd85, 8'd162, 8'd143, 8'd100, 8'd149, 8'd135, 8'd155, 8'd176, 8'd144, 8'd134, 8'd99, 8'd140, 8'd146, 8'd150, 8'd126, 8'd141, 8'd82, 8'd152, 8'd149, 8'd199, 8'd130, 8'd110, 8'd101, 8'd132, 8'd101, 8'd164, 8'd130, 8'd163, 8'd105, 8'd117, 8'd70, 8'd145, 8'd127, 8'd124, 8'd135, 8'd102, 8'd122, 8'd133, 8'd142, 8'd174, 8'd92, 8'd98, 8'd122, 8'd78, 8'd81, 8'd145, 8'd117, 8'd124, 8'd125, 8'd106, 8'd146, 8'd147, 8'd110, 8'd138, 8'd135, 8'd91, 8'd108, 8'd171, 8'd108, 8'd132, 8'd174, 8'd125, 8'd175, 8'd114, 8'd93, 8'd164, 8'd136, 8'd189, 8'd133, 8'd142, 8'd146, 8'd129, 8'd127, 8'd104, 8'd133, 8'd193, 8'd105, 8'd115, 8'd75, 8'd105, 8'd112, 8'd142, 8'd168, 8'd139, 8'd160, 8'd85, 8'd73, 8'd149, 8'd99, 8'd142, 8'd127, 8'd99, 8'd96, 8'd114, 8'd159, 8'd153, 8'd113, 8'd89, 8'd138, 8'd159, 8'd144, 8'd163, 8'd163, 8'd105, 8'd108, 8'd152, 8'd142, 8'd112, 8'd71, 8'd131, 8'd114, 8'd116, 8'd177, 8'd119, 8'd158, 8'd106, 8'd161, 8'd120, 8'd179, 8'd154, 8'd151, 8'd176, 8'd162, 8'd88, 8'd89, 8'd103, 8'd138, 8'd136, 8'd116, 8'd174, 8'd175, 8'd103, 8'd119, 8'd130, 8'd113, 8'd81, 8'd100, 8'd158, 8'd98, 8'd166, 8'd149, 8'd93, 8'd57, 8'd138, 8'd112, 8'd146, 8'd126, 8'd162, 8'd154, 8'd149, 8'd135, 8'd103, 8'd132, 8'd90, 8'd122, 8'd96, 8'd144, 8'd86, 8'd157, 8'd137, 8'd173, 8'd153, 8'd152, 8'd96, 8'd96, 8'd101, 8'd170, 8'd125, 8'd78, 8'd78, 8'd127, 8'd79, 8'd95, 8'd83, 8'd128, 8'd69, 8'd77, 8'd94, 8'd65, 8'd69, 8'd93, 8'd98, 8'd125, 8'd122, 8'd133, 8'd158, 8'd121, 8'd95, 8'd133, 8'd166, 8'd140, 8'd169, 8'd129, 8'd141, 8'd156, 8'd74, 8'd138, 8'd40, 8'd53, 8'd41, 8'd58, 8'd131, 8'd47, 8'd122, 8'd57, 8'd56, 8'd36, 8'd98, 8'd86, 8'd57, 8'd105, 8'd121, 8'd79, 8'd94, 8'd131, 8'd135, 8'd87, 8'd94, 8'd145, 8'd156, 8'd99, 8'd177, 8'd83, 8'd147, 8'd78, 8'd64, 8'd44, 8'd55, 8'd94, 8'd69, 8'd51, 8'd125, 8'd46, 8'd75, 8'd63, 8'd143, 8'd88, 8'd117, 8'd114, 8'd132, 8'd139, 8'd77, 8'd101, 8'd77, 8'd85, 8'd112, 8'd118, 8'd83, 8'd94, 8'd87, 8'd103, 8'd150, 8'd69, 8'd116, 8'd66, 8'd77, 8'd116, 8'd61, 8'd73, 8'd109, 8'd139, 8'd155, 8'd96, 8'd116, 8'd68, 8'd124, 8'd104, 8'd132, 8'd132, 8'd94, 8'd119, 8'd47, 8'd46, 8'd125, 8'd93, 8'd120, 8'd140, 8'd166, 8'd157, 8'd128, 8'd80, 8'd102, 8'd140, 8'd124, 8'd69, 8'd132, 8'd165, 8'd138, 8'd79, 8'd137, 8'd95, 8'd95, 8'd150, 8'd99, 8'd129, 8'd90, 8'd132, 8'd164, 8'd126, 8'd102, 8'd91, 8'd90, 8'd148, 8'd89, 8'd113, 8'd105, 8'd118, 8'd104, 8'd113, 8'd153, 8'd140, 8'd109, 8'd71, 8'd73, 8'd100, 8'd125, 8'd84, 8'd151, 8'd80, 8'd91, 8'd87, 8'd74, 8'd90, 8'd64, 8'd120, 8'd98, 8'd66, 8'd67, 8'd88, 8'd71, 8'd158, 8'd81, 8'd133, 8'd107, 8'd132, 8'd123, 8'd166, 8'd179, 8'd102, 8'd101, 8'd142, 8'd87, 8'd84, 8'd86, 8'd90, 8'd119, 8'd162, 8'd148, 8'd95, 8'd152, 8'd116, 8'd101, 8'd118, 8'd79, 8'd87, 8'd133, 8'd33, 8'd41, 8'd90, 8'd115, 8'd102, 8'd104, 8'd139, 8'd100, 8'd123, 8'd102, 8'd124, 8'd161, 8'd134, 8'd92, 8'd150, 8'd167, 8'd101, 8'd166, 8'd116, 8'd79, 8'd104, 8'd117, 8'd80, 8'd109, 8'd98, 8'd86, 8'd149, 8'd88, 8'd119, 8'd28, 8'd76, 8'd101, 8'd113, 8'd110, 8'd161, 8'd124, 8'd95, 8'd157, 8'd161, 8'd154, 8'd181, 8'd145, 8'd112, 8'd179, 8'd174, 8'd172, 8'd108, 8'd81, 8'd90, 8'd152, 8'd80, 8'd99, 8'd119, 8'd154, 8'd120, 8'd121, 8'd115, 8'd45, 8'd45, 8'd123, 8'd86, 8'd147, 8'd64, 8'd79, 8'd95, 8'd76, 8'd115, 8'd160, 8'd144, 8'd114, 8'd102, 8'd171, 8'd97, 8'd163, 8'd130, 8'd83, 8'd129, 8'd150, 8'd156, 8'd104, 8'd159, 8'd147, 8'd65, 8'd159, 8'd128, 8'd48, 8'd112, 8'd99, 8'd137, 8'd74, 8'd66, 8'd146, 8'd141, 8'd153, 8'd77, 8'd128, 8'd131, 8'd177, 8'd109, 8'd171, 8'd143, 8'd155, 8'd99, 8'd133, 8'd133, 8'd80, 8'd82, 8'd128, 8'd132, 8'd109, 8'd148, 8'd164, 8'd153, 8'd149, 8'd83, 8'd56, 8'd133, 8'd138, 8'd61, 8'd73, 8'd97, 8'd66, 8'd62, 8'd78, 8'd129, 8'd104, 8'd150, 8'd78, 8'd73, 8'd73, 8'd61, 8'd151, 8'd122, 8'd138, 8'd83, 8'd140, 8'd97, 8'd153, 8'd79, 8'd113, 8'd87, 8'd124, 8'd143, 8'd150, 8'd62, 8'd106, 8'd81, 8'd157, 8'd181, 8'd156, 8'd149, 8'd128, 8'd57, 8'd140, 8'd115, 8'd107, 8'd156, 8'd144, 8'd120, 8'd79, 8'd126, 8'd169, 8'd93, 8'd158, 8'd164, 8'd123, 8'd145, 8'd131, 8'd85, 8'd81, 8'd96, 8'd135, 8'd89, 8'd118, 8'd154, 8'd78, 8'd114, 8'd104, 8'd136, 8'd99, 8'd125, 8'd136, 8'd160, 8'd105, 8'd111, 8'd126, 8'd122, 8'd110, 8'd82, 8'd102, 8'd149, 8'd144, 8'd162})
) cell_0_79 (
    .clk(clk),
    .input_index(index_0_78_79),
    .input_value(value_0_78_79),
    .input_result(result_0_78_79),
    .input_enable(enable_0_78_79),
    .output_index(index_0_79_80),
    .output_value(value_0_79_80),
    .output_result(result_0_79_80),
    .output_enable(enable_0_79_80)
);

wire [10-1:0] index_0_80_81;
wire [`DATA_WIDTH-1:0] value_0_80_81;
wire [`DATA_WIDTH*4:0] result_0_80_81;
wire enable_0_80_81;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd103, 8'd93, 8'd168, 8'd156, 8'd83, 8'd146, 8'd122, 8'd122, 8'd145, 8'd104, 8'd123, 8'd121, 8'd105, 8'd84, 8'd104, 8'd116, 8'd102, 8'd85, 8'd93, 8'd96, 8'd150, 8'd106, 8'd103, 8'd111, 8'd131, 8'd88, 8'd79, 8'd130, 8'd95, 8'd106, 8'd158, 8'd74, 8'd148, 8'd123, 8'd79, 8'd88, 8'd128, 8'd74, 8'd42, 8'd84, 8'd74, 8'd72, 8'd97, 8'd94, 8'd117, 8'd38, 8'd73, 8'd72, 8'd104, 8'd82, 8'd141, 8'd115, 8'd140, 8'd100, 8'd140, 8'd155, 8'd102, 8'd117, 8'd139, 8'd80, 8'd74, 8'd55, 8'd85, 8'd71, 8'd86, 8'd89, 8'd44, 8'd59, 8'd53, 8'd116, 8'd58, 8'd139, 8'd56, 8'd76, 8'd71, 8'd58, 8'd69, 8'd71, 8'd120, 8'd110, 8'd158, 8'd88, 8'd139, 8'd166, 8'd79, 8'd128, 8'd106, 8'd115, 8'd139, 8'd106, 8'd129, 8'd111, 8'd95, 8'd111, 8'd104, 8'd121, 8'd83, 8'd135, 8'd121, 8'd133, 8'd101, 8'd147, 8'd148, 8'd104, 8'd88, 8'd145, 8'd130, 8'd181, 8'd126, 8'd152, 8'd149, 8'd149, 8'd86, 8'd177, 8'd103, 8'd97, 8'd83, 8'd139, 8'd120, 8'd83, 8'd171, 8'd102, 8'd105, 8'd152, 8'd102, 8'd113, 8'd87, 8'd144, 8'd148, 8'd126, 8'd112, 8'd80, 8'd175, 8'd159, 8'd107, 8'd172, 8'd172, 8'd181, 8'd149, 8'd151, 8'd82, 8'd127, 8'd68, 8'd110, 8'd74, 8'd153, 8'd120, 8'd162, 8'd125, 8'd148, 8'd169, 8'd161, 8'd93, 8'd127, 8'd156, 8'd90, 8'd158, 8'd142, 8'd110, 8'd91, 8'd102, 8'd82, 8'd89, 8'd160, 8'd98, 8'd178, 8'd115, 8'd125, 8'd124, 8'd154, 8'd69, 8'd127, 8'd72, 8'd112, 8'd77, 8'd80, 8'd118, 8'd92, 8'd115, 8'd133, 8'd144, 8'd93, 8'd110, 8'd109, 8'd170, 8'd101, 8'd171, 8'd105, 8'd117, 8'd162, 8'd91, 8'd157, 8'd136, 8'd176, 8'd173, 8'd138, 8'd143, 8'd87, 8'd154, 8'd107, 8'd112, 8'd73, 8'd166, 8'd166, 8'd97, 8'd99, 8'd94, 8'd102, 8'd93, 8'd138, 8'd132, 8'd164, 8'd100, 8'd178, 8'd125, 8'd138, 8'd166, 8'd147, 8'd103, 8'd165, 8'd118, 8'd132, 8'd141, 8'd126, 8'd129, 8'd79, 8'd139, 8'd91, 8'd85, 8'd124, 8'd133, 8'd104, 8'd174, 8'd170, 8'd188, 8'd144, 8'd143, 8'd115, 8'd169, 8'd79, 8'd100, 8'd171, 8'd155, 8'd166, 8'd87, 8'd106, 8'd119, 8'd130, 8'd180, 8'd110, 8'd76, 8'd139, 8'd86, 8'd76, 8'd175, 8'd143, 8'd176, 8'd164, 8'd108, 8'd149, 8'd180, 8'd185, 8'd147, 8'd127, 8'd133, 8'd130, 8'd158, 8'd74, 8'd151, 8'd75, 8'd162, 8'd171, 8'd85, 8'd98, 8'd101, 8'd109, 8'd153, 8'd110, 8'd122, 8'd88, 8'd116, 8'd80, 8'd137, 8'd161, 8'd154, 8'd99, 8'd160, 8'd121, 8'd130, 8'd133, 8'd164, 8'd90, 8'd85, 8'd152, 8'd59, 8'd67, 8'd96, 8'd84, 8'd99, 8'd172, 8'd113, 8'd117, 8'd158, 8'd96, 8'd182, 8'd121, 8'd134, 8'd86, 8'd90, 8'd105, 8'd106, 8'd164, 8'd143, 8'd156, 8'd168, 8'd117, 8'd162, 8'd142, 8'd71, 8'd73, 8'd78, 8'd165, 8'd67, 8'd123, 8'd98, 8'd149, 8'd111, 8'd94, 8'd96, 8'd122, 8'd111, 8'd104, 8'd109, 8'd107, 8'd171, 8'd67, 8'd88, 8'd97, 8'd110, 8'd181, 8'd111, 8'd114, 8'd94, 8'd95, 8'd135, 8'd133, 8'd102, 8'd117, 8'd128, 8'd149, 8'd118, 8'd130, 8'd130, 8'd98, 8'd163, 8'd175, 8'd175, 8'd126, 8'd145, 8'd85, 8'd123, 8'd150, 8'd149, 8'd132, 8'd91, 8'd116, 8'd172, 8'd154, 8'd207, 8'd125, 8'd165, 8'd98, 8'd120, 8'd158, 8'd92, 8'd143, 8'd98, 8'd92, 8'd94, 8'd166, 8'd199, 8'd106, 8'd167, 8'd140, 8'd150, 8'd152, 8'd107, 8'd106, 8'd101, 8'd103, 8'd93, 8'd94, 8'd148, 8'd75, 8'd106, 8'd218, 8'd182, 8'd111, 8'd145, 8'd99, 8'd127, 8'd120, 8'd134, 8'd108, 8'd159, 8'd177, 8'd153, 8'd173, 8'd135, 8'd125, 8'd96, 8'd104, 8'd173, 8'd73, 8'd134, 8'd93, 8'd90, 8'd97, 8'd124, 8'd81, 8'd128, 8'd137, 8'd103, 8'd164, 8'd182, 8'd168, 8'd118, 8'd115, 8'd75, 8'd96, 8'd88, 8'd69, 8'd125, 8'd81, 8'd96, 8'd155, 8'd143, 8'd162, 8'd88, 8'd139, 8'd69, 8'd65, 8'd132, 8'd45, 8'd70, 8'd103, 8'd114, 8'd108, 8'd165, 8'd125, 8'd81, 8'd79, 8'd141, 8'd84, 8'd135, 8'd87, 8'd83, 8'd85, 8'd112, 8'd145, 8'd148, 8'd115, 8'd130, 8'd158, 8'd115, 8'd81, 8'd97, 8'd126, 8'd83, 8'd94, 8'd45, 8'd129, 8'd84, 8'd130, 8'd156, 8'd145, 8'd88, 8'd61, 8'd145, 8'd87, 8'd149, 8'd117, 8'd118, 8'd112, 8'd158, 8'd87, 8'd109, 8'd82, 8'd115, 8'd99, 8'd106, 8'd88, 8'd45, 8'd104, 8'd90, 8'd110, 8'd111, 8'd53, 8'd81, 8'd91, 8'd171, 8'd125, 8'd118, 8'd149, 8'd119, 8'd62, 8'd78, 8'd56, 8'd87, 8'd69, 8'd77, 8'd117, 8'd92, 8'd107, 8'd114, 8'd114, 8'd95, 8'd117, 8'd61, 8'd53, 8'd78, 8'd139, 8'd70, 8'd129, 8'd80, 8'd69, 8'd100, 8'd152, 8'd161, 8'd104, 8'd120, 8'd130, 8'd153, 8'd118, 8'd113, 8'd81, 8'd133, 8'd122, 8'd68, 8'd146, 8'd83, 8'd148, 8'd63, 8'd82, 8'd146, 8'd96, 8'd74, 8'd88, 8'd65, 8'd130, 8'd64, 8'd79, 8'd73, 8'd79, 8'd112, 8'd179, 8'd93, 8'd149, 8'd98, 8'd112, 8'd152, 8'd139, 8'd49, 8'd99, 8'd67, 8'd95, 8'd111, 8'd118, 8'd144, 8'd68, 8'd139, 8'd88, 8'd91, 8'd115, 8'd109, 8'd111, 8'd146, 8'd133, 8'd59, 8'd109, 8'd74, 8'd91, 8'd119, 8'd189, 8'd172, 8'd160, 8'd83, 8'd80, 8'd123, 8'd83, 8'd99, 8'd148, 8'd177, 8'd125, 8'd138, 8'd161, 8'd106, 8'd92, 8'd164, 8'd80, 8'd104, 8'd62, 8'd129, 8'd137, 8'd127, 8'd153, 8'd134, 8'd79, 8'd78, 8'd121, 8'd114, 8'd144, 8'd110, 8'd136, 8'd92, 8'd119, 8'd122, 8'd121, 8'd75, 8'd159, 8'd160, 8'd98, 8'd178, 8'd168, 8'd108, 8'd139, 8'd169, 8'd112, 8'd121, 8'd101, 8'd153, 8'd135, 8'd161, 8'd121, 8'd116, 8'd140, 8'd152, 8'd138, 8'd151, 8'd102, 8'd150, 8'd122, 8'd128, 8'd105, 8'd77, 8'd158, 8'd120, 8'd104, 8'd105, 8'd128, 8'd175, 8'd107, 8'd149, 8'd147, 8'd118, 8'd121, 8'd164, 8'd185, 8'd96, 8'd112, 8'd107, 8'd125, 8'd127, 8'd151, 8'd110, 8'd105, 8'd129, 8'd108, 8'd101, 8'd143, 8'd94, 8'd71, 8'd160, 8'd85, 8'd142, 8'd171, 8'd174, 8'd99, 8'd165, 8'd167, 8'd142, 8'd136, 8'd179, 8'd171, 8'd109, 8'd184, 8'd206, 8'd146, 8'd126, 8'd178, 8'd175, 8'd171, 8'd179, 8'd123, 8'd101, 8'd132, 8'd82, 8'd138, 8'd124, 8'd121, 8'd129, 8'd91, 8'd121, 8'd173, 8'd95, 8'd172, 8'd114, 8'd105, 8'd145, 8'd126, 8'd164, 8'd136, 8'd131, 8'd153, 8'd166, 8'd142, 8'd200, 8'd186, 8'd158, 8'd160, 8'd111, 8'd151, 8'd130, 8'd138, 8'd159, 8'd133, 8'd135, 8'd143, 8'd89, 8'd167, 8'd164, 8'd94, 8'd114, 8'd145, 8'd157, 8'd132, 8'd93, 8'd110, 8'd174, 8'd90, 8'd145, 8'd92, 8'd159, 8'd151, 8'd169, 8'd158, 8'd166, 8'd91, 8'd166, 8'd168, 8'd109, 8'd153, 8'd142, 8'd132, 8'd147, 8'd110, 8'd113, 8'd155, 8'd75, 8'd168, 8'd154, 8'd109, 8'd112, 8'd132, 8'd129, 8'd136, 8'd132, 8'd118, 8'd118, 8'd131, 8'd122, 8'd160, 8'd157, 8'd72, 8'd99, 8'd166, 8'd102, 8'd131, 8'd82, 8'd86, 8'd162, 8'd157, 8'd119, 8'd161})
) cell_0_80 (
    .clk(clk),
    .input_index(index_0_79_80),
    .input_value(value_0_79_80),
    .input_result(result_0_79_80),
    .input_enable(enable_0_79_80),
    .output_index(index_0_80_81),
    .output_value(value_0_80_81),
    .output_result(result_0_80_81),
    .output_enable(enable_0_80_81)
);

wire [10-1:0] index_0_81_82;
wire [`DATA_WIDTH-1:0] value_0_81_82;
wire [`DATA_WIDTH*4:0] result_0_81_82;
wire enable_0_81_82;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd138, 8'd166, 8'd151, 8'd167, 8'd161, 8'd153, 8'd103, 8'd71, 8'd120, 8'd152, 8'd81, 8'd131, 8'd90, 8'd99, 8'd72, 8'd152, 8'd163, 8'd117, 8'd100, 8'd148, 8'd118, 8'd153, 8'd114, 8'd171, 8'd157, 8'd150, 8'd109, 8'd94, 8'd71, 8'd76, 8'd157, 8'd105, 8'd118, 8'd155, 8'd149, 8'd101, 8'd104, 8'd116, 8'd172, 8'd137, 8'd131, 8'd155, 8'd86, 8'd156, 8'd101, 8'd125, 8'd95, 8'd79, 8'd96, 8'd85, 8'd125, 8'd158, 8'd127, 8'd103, 8'd78, 8'd132, 8'd132, 8'd148, 8'd87, 8'd130, 8'd163, 8'd192, 8'd115, 8'd120, 8'd102, 8'd103, 8'd108, 8'd104, 8'd190, 8'd135, 8'd122, 8'd115, 8'd152, 8'd156, 8'd103, 8'd103, 8'd112, 8'd156, 8'd170, 8'd97, 8'd132, 8'd106, 8'd149, 8'd94, 8'd155, 8'd160, 8'd89, 8'd95, 8'd167, 8'd169, 8'd70, 8'd93, 8'd107, 8'd110, 8'd165, 8'd112, 8'd138, 8'd168, 8'd140, 8'd170, 8'd179, 8'd138, 8'd124, 8'd147, 8'd134, 8'd136, 8'd200, 8'd195, 8'd154, 8'd109, 8'd98, 8'd139, 8'd76, 8'd102, 8'd135, 8'd167, 8'd139, 8'd139, 8'd105, 8'd100, 8'd128, 8'd146, 8'd88, 8'd111, 8'd117, 8'd101, 8'd108, 8'd160, 8'd152, 8'd135, 8'd179, 8'd163, 8'd124, 8'd123, 8'd129, 8'd181, 8'd99, 8'd90, 8'd98, 8'd104, 8'd130, 8'd145, 8'd146, 8'd142, 8'd172, 8'd77, 8'd121, 8'd86, 8'd118, 8'd113, 8'd158, 8'd168, 8'd145, 8'd87, 8'd169, 8'd174, 8'd143, 8'd88, 8'd138, 8'd113, 8'd165, 8'd75, 8'd150, 8'd104, 8'd108, 8'd91, 8'd152, 8'd116, 8'd106, 8'd169, 8'd93, 8'd141, 8'd129, 8'd74, 8'd80, 8'd104, 8'd106, 8'd141, 8'd111, 8'd145, 8'd127, 8'd107, 8'd101, 8'd114, 8'd96, 8'd104, 8'd145, 8'd124, 8'd170, 8'd158, 8'd161, 8'd103, 8'd158, 8'd166, 8'd87, 8'd112, 8'd170, 8'd109, 8'd58, 8'd98, 8'd131, 8'd149, 8'd166, 8'd99, 8'd104, 8'd111, 8'd74, 8'd110, 8'd69, 8'd80, 8'd132, 8'd59, 8'd118, 8'd77, 8'd126, 8'd110, 8'd116, 8'd190, 8'd105, 8'd121, 8'd114, 8'd181, 8'd166, 8'd92, 8'd72, 8'd51, 8'd134, 8'd105, 8'd133, 8'd115, 8'd97, 8'd125, 8'd128, 8'd121, 8'd88, 8'd89, 8'd126, 8'd141, 8'd69, 8'd91, 8'd51, 8'd119, 8'd113, 8'd79, 8'd118, 8'd171, 8'd117, 8'd183, 8'd104, 8'd117, 8'd138, 8'd104, 8'd136, 8'd128, 8'd45, 8'd103, 8'd75, 8'd152, 8'd169, 8'd167, 8'd85, 8'd151, 8'd135, 8'd169, 8'd125, 8'd73, 8'd71, 8'd63, 8'd55, 8'd112, 8'd97, 8'd155, 8'd107, 8'd168, 8'd102, 8'd121, 8'd104, 8'd138, 8'd109, 8'd158, 8'd95, 8'd115, 8'd66, 8'd135, 8'd98, 8'd112, 8'd144, 8'd80, 8'd98, 8'd143, 8'd125, 8'd92, 8'd77, 8'd48, 8'd91, 8'd100, 8'd110, 8'd55, 8'd74, 8'd127, 8'd116, 8'd181, 8'd166, 8'd183, 8'd172, 8'd132, 8'd163, 8'd99, 8'd62, 8'd69, 8'd30, 8'd141, 8'd123, 8'd180, 8'd147, 8'd133, 8'd91, 8'd140, 8'd70, 8'd136, 8'd85, 8'd53, 8'd48, 8'd70, 8'd88, 8'd100, 8'd105, 8'd97, 8'd86, 8'd96, 8'd111, 8'd159, 8'd79, 8'd84, 8'd155, 8'd82, 8'd109, 8'd76, 8'd115, 8'd136, 8'd174, 8'd167, 8'd153, 8'd85, 8'd89, 8'd79, 8'd126, 8'd107, 8'd126, 8'd103, 8'd92, 8'd84, 8'd65, 8'd99, 8'd86, 8'd151, 8'd146, 8'd156, 8'd174, 8'd80, 8'd144, 8'd175, 8'd94, 8'd98, 8'd112, 8'd57, 8'd64, 8'd66, 8'd158, 8'd137, 8'd100, 8'd96, 8'd117, 8'd78, 8'd70, 8'd104, 8'd125, 8'd91, 8'd103, 8'd113, 8'd151, 8'd170, 8'd173, 8'd152, 8'd100, 8'd135, 8'd181, 8'd176, 8'd125, 8'd94, 8'd128, 8'd158, 8'd68, 8'd97, 8'd133, 8'd41, 8'd131, 8'd127, 8'd96, 8'd78, 8'd151, 8'd169, 8'd81, 8'd54, 8'd61, 8'd66, 8'd116, 8'd154, 8'd93, 8'd137, 8'd76, 8'd83, 8'd164, 8'd93, 8'd115, 8'd137, 8'd86, 8'd95, 8'd109, 8'd76, 8'd91, 8'd155, 8'd114, 8'd85, 8'd39, 8'd103, 8'd52, 8'd109, 8'd159, 8'd103, 8'd75, 8'd106, 8'd73, 8'd128, 8'd155, 8'd181, 8'd128, 8'd98, 8'd91, 8'd134, 8'd97, 8'd101, 8'd153, 8'd125, 8'd153, 8'd81, 8'd161, 8'd69, 8'd155, 8'd107, 8'd125, 8'd171, 8'd80, 8'd110, 8'd55, 8'd66, 8'd132, 8'd98, 8'd85, 8'd115, 8'd148, 8'd148, 8'd184, 8'd120, 8'd170, 8'd104, 8'd66, 8'd122, 8'd158, 8'd98, 8'd110, 8'd98, 8'd84, 8'd133, 8'd148, 8'd97, 8'd121, 8'd175, 8'd183, 8'd135, 8'd148, 8'd162, 8'd103, 8'd172, 8'd105, 8'd121, 8'd159, 8'd80, 8'd132, 8'd99, 8'd168, 8'd132, 8'd93, 8'd147, 8'd73, 8'd98, 8'd118, 8'd93, 8'd133, 8'd114, 8'd143, 8'd81, 8'd95, 8'd163, 8'd142, 8'd144, 8'd152, 8'd129, 8'd115, 8'd146, 8'd102, 8'd96, 8'd123, 8'd144, 8'd140, 8'd179, 8'd166, 8'd127, 8'd82, 8'd96, 8'd150, 8'd110, 8'd99, 8'd118, 8'd119, 8'd148, 8'd86, 8'd127, 8'd82, 8'd145, 8'd83, 8'd83, 8'd106, 8'd135, 8'd138, 8'd129, 8'd181, 8'd120, 8'd84, 8'd131, 8'd127, 8'd183, 8'd167, 8'd122, 8'd136, 8'd110, 8'd176, 8'd146, 8'd102, 8'd135, 8'd128, 8'd133, 8'd100, 8'd84, 8'd83, 8'd72, 8'd131, 8'd152, 8'd89, 8'd102, 8'd141, 8'd96, 8'd103, 8'd128, 8'd152, 8'd105, 8'd92, 8'd174, 8'd151, 8'd120, 8'd136, 8'd135, 8'd157, 8'd136, 8'd178, 8'd84, 8'd158, 8'd159, 8'd131, 8'd146, 8'd69, 8'd76, 8'd68, 8'd126, 8'd99, 8'd108, 8'd142, 8'd142, 8'd149, 8'd113, 8'd130, 8'd98, 8'd127, 8'd107, 8'd126, 8'd138, 8'd118, 8'd180, 8'd106, 8'd145, 8'd109, 8'd117, 8'd130, 8'd164, 8'd127, 8'd120, 8'd125, 8'd133, 8'd118, 8'd129, 8'd64, 8'd88, 8'd129, 8'd110, 8'd93, 8'd110, 8'd70, 8'd99, 8'd80, 8'd114, 8'd106, 8'd141, 8'd84, 8'd110, 8'd160, 8'd144, 8'd148, 8'd78, 8'd63, 8'd92, 8'd113, 8'd109, 8'd137, 8'd127, 8'd144, 8'd91, 8'd156, 8'd130, 8'd58, 8'd143, 8'd77, 8'd122, 8'd79, 8'd130, 8'd151, 8'd83, 8'd89, 8'd76, 8'd104, 8'd124, 8'd78, 8'd143, 8'd121, 8'd83, 8'd148, 8'd137, 8'd135, 8'd126, 8'd115, 8'd69, 8'd109, 8'd153, 8'd60, 8'd145, 8'd142, 8'd62, 8'd77, 8'd131, 8'd162, 8'd86, 8'd91, 8'd112, 8'd70, 8'd137, 8'd71, 8'd79, 8'd144, 8'd84, 8'd84, 8'd134, 8'd150, 8'd78, 8'd140, 8'd51, 8'd67, 8'd148, 8'd81, 8'd116, 8'd48, 8'd62, 8'd125, 8'd77, 8'd52, 8'd48, 8'd95, 8'd92, 8'd163, 8'd75, 8'd142, 8'd99, 8'd167, 8'd95, 8'd127, 8'd106, 8'd58, 8'd93, 8'd59, 8'd64, 8'd73, 8'd97, 8'd63, 8'd125, 8'd34, 8'd57, 8'd19, 8'd33, 8'd43, 8'd88, 8'd32, 8'd81, 8'd145, 8'd63, 8'd130, 8'd88, 8'd106, 8'd114, 8'd93, 8'd97, 8'd100, 8'd99, 8'd90, 8'd170, 8'd97, 8'd124, 8'd130, 8'd122, 8'd111, 8'd85, 8'd107, 8'd114, 8'd85, 8'd58, 8'd112, 8'd113, 8'd102, 8'd64, 8'd90, 8'd111, 8'd140, 8'd129, 8'd142, 8'd143, 8'd126, 8'd167, 8'd78, 8'd105, 8'd162, 8'd160, 8'd116, 8'd103, 8'd70, 8'd163, 8'd162, 8'd113, 8'd123, 8'd125, 8'd154, 8'd100, 8'd79, 8'd131, 8'd81, 8'd70, 8'd119, 8'd95, 8'd138, 8'd82, 8'd101, 8'd95, 8'd126, 8'd75, 8'd95, 8'd152, 8'd136, 8'd98})
) cell_0_81 (
    .clk(clk),
    .input_index(index_0_80_81),
    .input_value(value_0_80_81),
    .input_result(result_0_80_81),
    .input_enable(enable_0_80_81),
    .output_index(index_0_81_82),
    .output_value(value_0_81_82),
    .output_result(result_0_81_82),
    .output_enable(enable_0_81_82)
);

wire [10-1:0] index_0_82_83;
wire [`DATA_WIDTH-1:0] value_0_82_83;
wire [`DATA_WIDTH*4:0] result_0_82_83;
wire enable_0_82_83;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd159, 8'd112, 8'd113, 8'd72, 8'd82, 8'd96, 8'd101, 8'd168, 8'd173, 8'd109, 8'd123, 8'd166, 8'd165, 8'd184, 8'd131, 8'd80, 8'd159, 8'd149, 8'd145, 8'd103, 8'd142, 8'd127, 8'd99, 8'd132, 8'd119, 8'd99, 8'd168, 8'd76, 8'd96, 8'd118, 8'd82, 8'd142, 8'd142, 8'd107, 8'd133, 8'd85, 8'd112, 8'd161, 8'd152, 8'd80, 8'd99, 8'd98, 8'd115, 8'd109, 8'd115, 8'd96, 8'd71, 8'd72, 8'd107, 8'd86, 8'd72, 8'd88, 8'd108, 8'd86, 8'd145, 8'd134, 8'd146, 8'd94, 8'd64, 8'd146, 8'd104, 8'd82, 8'd138, 8'd57, 8'd159, 8'd58, 8'd88, 8'd53, 8'd74, 8'd105, 8'd156, 8'd72, 8'd81, 8'd165, 8'd121, 8'd84, 8'd150, 8'd157, 8'd88, 8'd130, 8'd119, 8'd157, 8'd110, 8'd98, 8'd133, 8'd154, 8'd70, 8'd71, 8'd62, 8'd39, 8'd115, 8'd126, 8'd136, 8'd74, 8'd160, 8'd115, 8'd159, 8'd164, 8'd157, 8'd168, 8'd120, 8'd129, 8'd77, 8'd159, 8'd175, 8'd109, 8'd151, 8'd93, 8'd159, 8'd72, 8'd79, 8'd110, 8'd128, 8'd112, 8'd140, 8'd59, 8'd99, 8'd133, 8'd115, 8'd68, 8'd95, 8'd160, 8'd162, 8'd128, 8'd156, 8'd188, 8'd146, 8'd95, 8'd81, 8'd110, 8'd143, 8'd148, 8'd108, 8'd77, 8'd153, 8'd106, 8'd98, 8'd100, 8'd132, 8'd82, 8'd79, 8'd167, 8'd131, 8'd42, 8'd52, 8'd136, 8'd85, 8'd112, 8'd96, 8'd137, 8'd127, 8'd81, 8'd145, 8'd95, 8'd125, 8'd117, 8'd142, 8'd104, 8'd154, 8'd97, 8'd65, 8'd118, 8'd122, 8'd124, 8'd110, 8'd147, 8'd125, 8'd128, 8'd105, 8'd139, 8'd81, 8'd102, 8'd104, 8'd99, 8'd122, 8'd100, 8'd67, 8'd59, 8'd129, 8'd160, 8'd149, 8'd152, 8'd111, 8'd141, 8'd169, 8'd115, 8'd104, 8'd73, 8'd106, 8'd67, 8'd99, 8'd139, 8'd75, 8'd103, 8'd91, 8'd129, 8'd129, 8'd104, 8'd42, 8'd113, 8'd49, 8'd101, 8'd144, 8'd150, 8'd143, 8'd68, 8'd121, 8'd158, 8'd134, 8'd127, 8'd156, 8'd115, 8'd106, 8'd86, 8'd84, 8'd90, 8'd109, 8'd133, 8'd82, 8'd139, 8'd137, 8'd159, 8'd78, 8'd164, 8'd150, 8'd129, 8'd101, 8'd74, 8'd78, 8'd115, 8'd152, 8'd153, 8'd130, 8'd151, 8'd126, 8'd101, 8'd97, 8'd62, 8'd92, 8'd109, 8'd115, 8'd119, 8'd111, 8'd140, 8'd143, 8'd70, 8'd108, 8'd85, 8'd134, 8'd154, 8'd166, 8'd152, 8'd124, 8'd77, 8'd126, 8'd101, 8'd109, 8'd132, 8'd144, 8'd160, 8'd131, 8'd162, 8'd71, 8'd84, 8'd146, 8'd115, 8'd90, 8'd110, 8'd136, 8'd132, 8'd121, 8'd143, 8'd143, 8'd137, 8'd74, 8'd133, 8'd119, 8'd160, 8'd144, 8'd168, 8'd82, 8'd104, 8'd69, 8'd118, 8'd147, 8'd161, 8'd78, 8'd165, 8'd154, 8'd91, 8'd96, 8'd131, 8'd146, 8'd112, 8'd78, 8'd92, 8'd83, 8'd142, 8'd107, 8'd165, 8'd155, 8'd94, 8'd107, 8'd143, 8'd74, 8'd90, 8'd129, 8'd169, 8'd107, 8'd61, 8'd56, 8'd134, 8'd85, 8'd91, 8'd137, 8'd103, 8'd178, 8'd135, 8'd107, 8'd119, 8'd124, 8'd135, 8'd49, 8'd109, 8'd133, 8'd146, 8'd199, 8'd115, 8'd194, 8'd161, 8'd75, 8'd101, 8'd123, 8'd87, 8'd82, 8'd118, 8'd93, 8'd122, 8'd81, 8'd97, 8'd146, 8'd136, 8'd106, 8'd103, 8'd175, 8'd142, 8'd94, 8'd77, 8'd114, 8'd94, 8'd51, 8'd148, 8'd142, 8'd91, 8'd101, 8'd186, 8'd191, 8'd164, 8'd113, 8'd118, 8'd86, 8'd183, 8'd119, 8'd110, 8'd109, 8'd77, 8'd140, 8'd155, 8'd100, 8'd105, 8'd140, 8'd107, 8'd96, 8'd119, 8'd172, 8'd146, 8'd137, 8'd109, 8'd56, 8'd94, 8'd116, 8'd162, 8'd179, 8'd158, 8'd117, 8'd145, 8'd157, 8'd129, 8'd122, 8'd167, 8'd155, 8'd131, 8'd75, 8'd105, 8'd100, 8'd118, 8'd157, 8'd108, 8'd92, 8'd107, 8'd129, 8'd147, 8'd131, 8'd130, 8'd84, 8'd135, 8'd113, 8'd102, 8'd182, 8'd105, 8'd191, 8'd130, 8'd181, 8'd184, 8'd162, 8'd92, 8'd169, 8'd166, 8'd167, 8'd90, 8'd82, 8'd71, 8'd151, 8'd127, 8'd144, 8'd158, 8'd105, 8'd122, 8'd117, 8'd128, 8'd137, 8'd81, 8'd120, 8'd64, 8'd87, 8'd113, 8'd149, 8'd149, 8'd113, 8'd153, 8'd140, 8'd105, 8'd93, 8'd107, 8'd151, 8'd101, 8'd177, 8'd89, 8'd120, 8'd53, 8'd46, 8'd150, 8'd115, 8'd113, 8'd124, 8'd173, 8'd162, 8'd155, 8'd174, 8'd94, 8'd146, 8'd116, 8'd108, 8'd106, 8'd135, 8'd153, 8'd164, 8'd111, 8'd175, 8'd120, 8'd126, 8'd87, 8'd176, 8'd147, 8'd132, 8'd79, 8'd145, 8'd34, 8'd7, 8'd79, 8'd157, 8'd109, 8'd126, 8'd149, 8'd105, 8'd181, 8'd137, 8'd83, 8'd88, 8'd101, 8'd153, 8'd166, 8'd165, 8'd95, 8'd144, 8'd140, 8'd138, 8'd161, 8'd150, 8'd91, 8'd111, 8'd140, 8'd163, 8'd159, 8'd72, 8'd81, 8'd36, 8'd67, 8'd163, 8'd122, 8'd146, 8'd130, 8'd96, 8'd107, 8'd106, 8'd81, 8'd142, 8'd105, 8'd71, 8'd114, 8'd129, 8'd156, 8'd59, 8'd84, 8'd132, 8'd129, 8'd91, 8'd151, 8'd150, 8'd90, 8'd109, 8'd106, 8'd151, 8'd62, 8'd51, 8'd87, 8'd92, 8'd140, 8'd153, 8'd90, 8'd94, 8'd175, 8'd130, 8'd155, 8'd105, 8'd128, 8'd128, 8'd72, 8'd91, 8'd102, 8'd106, 8'd69, 8'd144, 8'd167, 8'd140, 8'd122, 8'd96, 8'd154, 8'd127, 8'd165, 8'd78, 8'd61, 8'd81, 8'd152, 8'd91, 8'd81, 8'd141, 8'd128, 8'd161, 8'd117, 8'd95, 8'd131, 8'd125, 8'd105, 8'd77, 8'd70, 8'd107, 8'd79, 8'd85, 8'd75, 8'd131, 8'd164, 8'd110, 8'd123, 8'd100, 8'd136, 8'd98, 8'd137, 8'd87, 8'd119, 8'd104, 8'd110, 8'd111, 8'd137, 8'd157, 8'd88, 8'd154, 8'd82, 8'd130, 8'd149, 8'd93, 8'd118, 8'd159, 8'd122, 8'd83, 8'd158, 8'd75, 8'd144, 8'd147, 8'd132, 8'd119, 8'd136, 8'd157, 8'd132, 8'd118, 8'd131, 8'd130, 8'd155, 8'd104, 8'd137, 8'd166, 8'd126, 8'd89, 8'd150, 8'd127, 8'd136, 8'd80, 8'd116, 8'd66, 8'd146, 8'd81, 8'd121, 8'd119, 8'd138, 8'd115, 8'd109, 8'd100, 8'd96, 8'd127, 8'd85, 8'd161, 8'd78, 8'd87, 8'd147, 8'd110, 8'd121, 8'd83, 8'd142, 8'd117, 8'd113, 8'd81, 8'd98, 8'd152, 8'd119, 8'd150, 8'd97, 8'd131, 8'd145, 8'd104, 8'd111, 8'd133, 8'd80, 8'd97, 8'd100, 8'd128, 8'd158, 8'd103, 8'd130, 8'd131, 8'd148, 8'd93, 8'd71, 8'd101, 8'd122, 8'd153, 8'd114, 8'd123, 8'd163, 8'd123, 8'd108, 8'd85, 8'd125, 8'd146, 8'd85, 8'd135, 8'd157, 8'd148, 8'd99, 8'd150, 8'd115, 8'd106, 8'd96, 8'd140, 8'd153, 8'd124, 8'd118, 8'd122, 8'd148, 8'd156, 8'd116, 8'd158, 8'd162, 8'd134, 8'd163, 8'd172, 8'd157, 8'd172, 8'd152, 8'd115, 8'd166, 8'd148, 8'd118, 8'd128, 8'd150, 8'd166, 8'd159, 8'd135, 8'd107, 8'd115, 8'd147, 8'd121, 8'd173, 8'd101, 8'd137, 8'd172, 8'd76, 8'd113, 8'd82, 8'd148, 8'd109, 8'd87, 8'd124, 8'd115, 8'd120, 8'd159, 8'd155, 8'd138, 8'd175, 8'd139, 8'd126, 8'd168, 8'd154, 8'd131, 8'd121, 8'd182, 8'd155, 8'd128, 8'd146, 8'd142, 8'd109, 8'd133, 8'd156, 8'd70, 8'd152, 8'd81, 8'd103, 8'd140, 8'd120, 8'd115, 8'd95, 8'd78, 8'd70, 8'd83, 8'd164, 8'd95, 8'd118, 8'd74, 8'd138, 8'd137, 8'd113, 8'd147, 8'd113, 8'd75, 8'd140, 8'd116, 8'd113, 8'd77, 8'd99, 8'd139, 8'd97, 8'd87, 8'd80, 8'd120, 8'd73})
) cell_0_82 (
    .clk(clk),
    .input_index(index_0_81_82),
    .input_value(value_0_81_82),
    .input_result(result_0_81_82),
    .input_enable(enable_0_81_82),
    .output_index(index_0_82_83),
    .output_value(value_0_82_83),
    .output_result(result_0_82_83),
    .output_enable(enable_0_82_83)
);

wire [10-1:0] index_0_83_84;
wire [`DATA_WIDTH-1:0] value_0_83_84;
wire [`DATA_WIDTH*4:0] result_0_83_84;
wire enable_0_83_84;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd103, 8'd103, 8'd144, 8'd99, 8'd155, 8'd159, 8'd134, 8'd174, 8'd87, 8'd95, 8'd106, 8'd177, 8'd127, 8'd131, 8'd90, 8'd83, 8'd119, 8'd90, 8'd131, 8'd112, 8'd176, 8'd89, 8'd74, 8'd98, 8'd91, 8'd73, 8'd165, 8'd168, 8'd106, 8'd88, 8'd164, 8'd160, 8'd138, 8'd175, 8'd134, 8'd152, 8'd166, 8'd171, 8'd122, 8'd166, 8'd124, 8'd153, 8'd201, 8'd212, 8'd174, 8'd159, 8'd166, 8'd175, 8'd104, 8'd181, 8'd131, 8'd117, 8'd112, 8'd138, 8'd139, 8'd168, 8'd70, 8'd101, 8'd162, 8'd93, 8'd172, 8'd117, 8'd99, 8'd136, 8'd117, 8'd158, 8'd132, 8'd148, 8'd119, 8'd138, 8'd109, 8'd103, 8'd122, 8'd127, 8'd169, 8'd101, 8'd106, 8'd156, 8'd106, 8'd144, 8'd129, 8'd125, 8'd164, 8'd75, 8'd98, 8'd92, 8'd105, 8'd104, 8'd129, 8'd170, 8'd75, 8'd171, 8'd123, 8'd150, 8'd104, 8'd63, 8'd96, 8'd142, 8'd73, 8'd157, 8'd105, 8'd106, 8'd118, 8'd134, 8'd72, 8'd99, 8'd119, 8'd66, 8'd64, 8'd68, 8'd77, 8'd126, 8'd74, 8'd135, 8'd68, 8'd106, 8'd90, 8'd137, 8'd76, 8'd76, 8'd68, 8'd91, 8'd116, 8'd101, 8'd122, 8'd79, 8'd136, 8'd69, 8'd114, 8'd73, 8'd73, 8'd157, 8'd121, 8'd103, 8'd97, 8'd71, 8'd81, 8'd133, 8'd80, 8'd113, 8'd146, 8'd75, 8'd146, 8'd119, 8'd91, 8'd74, 8'd123, 8'd116, 8'd136, 8'd61, 8'd89, 8'd79, 8'd113, 8'd163, 8'd123, 8'd152, 8'd84, 8'd155, 8'd157, 8'd152, 8'd106, 8'd94, 8'd92, 8'd138, 8'd124, 8'd130, 8'd142, 8'd111, 8'd100, 8'd138, 8'd94, 8'd99, 8'd70, 8'd131, 8'd135, 8'd115, 8'd79, 8'd105, 8'd144, 8'd119, 8'd99, 8'd119, 8'd99, 8'd164, 8'd103, 8'd98, 8'd115, 8'd106, 8'd151, 8'd85, 8'd109, 8'd82, 8'd127, 8'd117, 8'd166, 8'd85, 8'd153, 8'd107, 8'd120, 8'd85, 8'd91, 8'd70, 8'd72, 8'd145, 8'd89, 8'd101, 8'd112, 8'd101, 8'd82, 8'd143, 8'd169, 8'd161, 8'd121, 8'd134, 8'd130, 8'd143, 8'd65, 8'd83, 8'd152, 8'd121, 8'd110, 8'd134, 8'd155, 8'd148, 8'd81, 8'd90, 8'd76, 8'd83, 8'd123, 8'd116, 8'd128, 8'd140, 8'd134, 8'd135, 8'd81, 8'd153, 8'd150, 8'd152, 8'd104, 8'd117, 8'd138, 8'd109, 8'd172, 8'd89, 8'd99, 8'd67, 8'd64, 8'd95, 8'd111, 8'd98, 8'd115, 8'd105, 8'd139, 8'd151, 8'd78, 8'd148, 8'd64, 8'd161, 8'd140, 8'd148, 8'd84, 8'd153, 8'd94, 8'd81, 8'd61, 8'd93, 8'd68, 8'd97, 8'd101, 8'd147, 8'd145, 8'd126, 8'd103, 8'd145, 8'd109, 8'd63, 8'd135, 8'd108, 8'd156, 8'd180, 8'd150, 8'd83, 8'd76, 8'd58, 8'd96, 8'd79, 8'd153, 8'd111, 8'd92, 8'd99, 8'd87, 8'd151, 8'd120, 8'd65, 8'd75, 8'd113, 8'd155, 8'd139, 8'd127, 8'd160, 8'd86, 8'd146, 8'd110, 8'd141, 8'd128, 8'd124, 8'd129, 8'd86, 8'd73, 8'd59, 8'd119, 8'd68, 8'd140, 8'd93, 8'd79, 8'd98, 8'd109, 8'd142, 8'd64, 8'd94, 8'd108, 8'd65, 8'd91, 8'd127, 8'd80, 8'd168, 8'd102, 8'd157, 8'd162, 8'd91, 8'd152, 8'd82, 8'd85, 8'd57, 8'd85, 8'd141, 8'd96, 8'd55, 8'd71, 8'd102, 8'd166, 8'd141, 8'd150, 8'd123, 8'd137, 8'd145, 8'd134, 8'd57, 8'd108, 8'd120, 8'd84, 8'd96, 8'd145, 8'd160, 8'd100, 8'd87, 8'd77, 8'd87, 8'd112, 8'd67, 8'd80, 8'd98, 8'd105, 8'd120, 8'd157, 8'd119, 8'd131, 8'd145, 8'd123, 8'd121, 8'd128, 8'd142, 8'd60, 8'd70, 8'd130, 8'd111, 8'd95, 8'd143, 8'd98, 8'd125, 8'd102, 8'd112, 8'd163, 8'd139, 8'd171, 8'd173, 8'd135, 8'd97, 8'd117, 8'd82, 8'd113, 8'd116, 8'd131, 8'd92, 8'd133, 8'd86, 8'd112, 8'd95, 8'd118, 8'd86, 8'd107, 8'd149, 8'd115, 8'd88, 8'd150, 8'd146, 8'd128, 8'd142, 8'd73, 8'd153, 8'd110, 8'd110, 8'd87, 8'd124, 8'd153, 8'd134, 8'd110, 8'd97, 8'd80, 8'd131, 8'd97, 8'd119, 8'd124, 8'd139, 8'd161, 8'd168, 8'd94, 8'd165, 8'd97, 8'd115, 8'd66, 8'd121, 8'd121, 8'd102, 8'd123, 8'd101, 8'd118, 8'd154, 8'd166, 8'd126, 8'd174, 8'd112, 8'd106, 8'd141, 8'd133, 8'd92, 8'd175, 8'd69, 8'd98, 8'd49, 8'd42, 8'd160, 8'd162, 8'd87, 8'd168, 8'd138, 8'd110, 8'd129, 8'd88, 8'd123, 8'd85, 8'd119, 8'd123, 8'd135, 8'd140, 8'd161, 8'd101, 8'd123, 8'd148, 8'd129, 8'd140, 8'd81, 8'd144, 8'd174, 8'd177, 8'd117, 8'd140, 8'd107, 8'd84, 8'd146, 8'd130, 8'd140, 8'd102, 8'd69, 8'd59, 8'd106, 8'd122, 8'd110, 8'd103, 8'd158, 8'd159, 8'd161, 8'd83, 8'd109, 8'd141, 8'd174, 8'd168, 8'd150, 8'd127, 8'd157, 8'd117, 8'd171, 8'd103, 8'd129, 8'd140, 8'd96, 8'd133, 8'd80, 8'd138, 8'd91, 8'd145, 8'd81, 8'd154, 8'd114, 8'd145, 8'd124, 8'd86, 8'd182, 8'd163, 8'd163, 8'd117, 8'd91, 8'd137, 8'd94, 8'd115, 8'd97, 8'd148, 8'd101, 8'd100, 8'd67, 8'd95, 8'd90, 8'd94, 8'd137, 8'd70, 8'd140, 8'd99, 8'd110, 8'd113, 8'd70, 8'd123, 8'd122, 8'd150, 8'd155, 8'd162, 8'd160, 8'd137, 8'd162, 8'd155, 8'd77, 8'd62, 8'd68, 8'd78, 8'd110, 8'd131, 8'd53, 8'd73, 8'd98, 8'd75, 8'd161, 8'd136, 8'd145, 8'd136, 8'd148, 8'd154, 8'd161, 8'd73, 8'd78, 8'd132, 8'd151, 8'd130, 8'd115, 8'd145, 8'd109, 8'd122, 8'd79, 8'd82, 8'd123, 8'd134, 8'd147, 8'd62, 8'd90, 8'd104, 8'd84, 8'd124, 8'd85, 8'd101, 8'd155, 8'd109, 8'd123, 8'd120, 8'd115, 8'd118, 8'd102, 8'd175, 8'd91, 8'd168, 8'd109, 8'd107, 8'd132, 8'd110, 8'd102, 8'd171, 8'd104, 8'd164, 8'd60, 8'd53, 8'd127, 8'd110, 8'd135, 8'd122, 8'd47, 8'd118, 8'd157, 8'd123, 8'd166, 8'd132, 8'd133, 8'd124, 8'd161, 8'd106, 8'd119, 8'd100, 8'd106, 8'd130, 8'd67, 8'd70, 8'd121, 8'd89, 8'd160, 8'd148, 8'd93, 8'd96, 8'd140, 8'd115, 8'd141, 8'd57, 8'd144, 8'd118, 8'd73, 8'd66, 8'd72, 8'd76, 8'd151, 8'd147, 8'd90, 8'd101, 8'd144, 8'd160, 8'd116, 8'd118, 8'd151, 8'd84, 8'd96, 8'd144, 8'd96, 8'd122, 8'd65, 8'd88, 8'd132, 8'd58, 8'd91, 8'd140, 8'd149, 8'd143, 8'd128, 8'd112, 8'd115, 8'd79, 8'd81, 8'd156, 8'd71, 8'd104, 8'd81, 8'd155, 8'd150, 8'd187, 8'd115, 8'd154, 8'd134, 8'd116, 8'd92, 8'd151, 8'd139, 8'd121, 8'd108, 8'd100, 8'd138, 8'd123, 8'd107, 8'd157, 8'd80, 8'd90, 8'd115, 8'd127, 8'd170, 8'd94, 8'd141, 8'd138, 8'd117, 8'd153, 8'd103, 8'd154, 8'd140, 8'd165, 8'd167, 8'd155, 8'd168, 8'd137, 8'd173, 8'd171, 8'd142, 8'd112, 8'd104, 8'd163, 8'd97, 8'd143, 8'd109, 8'd105, 8'd190, 8'd183, 8'd110, 8'd108, 8'd137, 8'd122, 8'd110, 8'd146, 8'd136, 8'd98, 8'd80, 8'd142, 8'd98, 8'd93, 8'd88, 8'd104, 8'd102, 8'd88, 8'd183, 8'd176, 8'd148, 8'd177, 8'd80, 8'd166, 8'd139, 8'd108, 8'd93, 8'd112, 8'd167, 8'd113, 8'd124, 8'd128, 8'd136, 8'd77, 8'd80, 8'd91, 8'd138, 8'd139, 8'd166, 8'd113, 8'd152, 8'd78, 8'd83, 8'd73, 8'd139, 8'd161, 8'd137, 8'd146, 8'd91, 8'd100, 8'd130, 8'd147, 8'd121, 8'd85, 8'd165, 8'd122, 8'd159, 8'd83, 8'd95, 8'd139, 8'd94, 8'd154, 8'd145, 8'd116, 8'd97})
) cell_0_83 (
    .clk(clk),
    .input_index(index_0_82_83),
    .input_value(value_0_82_83),
    .input_result(result_0_82_83),
    .input_enable(enable_0_82_83),
    .output_index(index_0_83_84),
    .output_value(value_0_83_84),
    .output_result(result_0_83_84),
    .output_enable(enable_0_83_84)
);

wire [10-1:0] index_0_84_85;
wire [`DATA_WIDTH-1:0] value_0_84_85;
wire [`DATA_WIDTH*4:0] result_0_84_85;
wire enable_0_84_85;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd111, 8'd95, 8'd76, 8'd79, 8'd109, 8'd73, 8'd77, 8'd155, 8'd70, 8'd124, 8'd121, 8'd108, 8'd61, 8'd137, 8'd69, 8'd114, 8'd131, 8'd141, 8'd103, 8'd154, 8'd120, 8'd128, 8'd144, 8'd153, 8'd85, 8'd121, 8'd126, 8'd143, 8'd81, 8'd112, 8'd161, 8'd135, 8'd107, 8'd119, 8'd94, 8'd86, 8'd65, 8'd63, 8'd90, 8'd133, 8'd143, 8'd128, 8'd139, 8'd100, 8'd136, 8'd78, 8'd119, 8'd110, 8'd165, 8'd152, 8'd115, 8'd91, 8'd86, 8'd159, 8'd105, 8'd137, 8'd95, 8'd88, 8'd94, 8'd98, 8'd99, 8'd97, 8'd139, 8'd102, 8'd155, 8'd64, 8'd127, 8'd65, 8'd95, 8'd89, 8'd107, 8'd33, 8'd121, 8'd48, 8'd110, 8'd64, 8'd76, 8'd112, 8'd89, 8'd102, 8'd153, 8'd88, 8'd94, 8'd150, 8'd146, 8'd88, 8'd144, 8'd152, 8'd112, 8'd98, 8'd122, 8'd134, 8'd73, 8'd73, 8'd46, 8'd98, 8'd53, 8'd95, 8'd27, 8'd117, 8'd118, 8'd121, 8'd96, 8'd117, 8'd110, 8'd110, 8'd52, 8'd49, 8'd38, 8'd157, 8'd127, 8'd157, 8'd94, 8'd111, 8'd132, 8'd145, 8'd110, 8'd119, 8'd184, 8'd162, 8'd117, 8'd101, 8'd113, 8'd92, 8'd120, 8'd89, 8'd64, 8'd75, 8'd60, 8'd94, 8'd98, 8'd79, 8'd75, 8'd54, 8'd109, 8'd113, 8'd124, 8'd104, 8'd133, 8'd88, 8'd148, 8'd161, 8'd80, 8'd179, 8'd102, 8'd146, 8'd89, 8'd158, 8'd127, 8'd90, 8'd66, 8'd164, 8'd106, 8'd113, 8'd78, 8'd156, 8'd99, 8'd151, 8'd96, 8'd79, 8'd95, 8'd75, 8'd67, 8'd87, 8'd156, 8'd82, 8'd104, 8'd89, 8'd139, 8'd134, 8'd158, 8'd149, 8'd179, 8'd153, 8'd173, 8'd175, 8'd112, 8'd180, 8'd100, 8'd144, 8'd164, 8'd91, 8'd159, 8'd176, 8'd92, 8'd152, 8'd111, 8'd81, 8'd89, 8'd154, 8'd160, 8'd125, 8'd129, 8'd100, 8'd121, 8'd149, 8'd140, 8'd114, 8'd137, 8'd173, 8'd117, 8'd135, 8'd123, 8'd183, 8'd185, 8'd102, 8'd169, 8'd112, 8'd165, 8'd181, 8'd164, 8'd178, 8'd194, 8'd202, 8'd154, 8'd164, 8'd116, 8'd81, 8'd118, 8'd56, 8'd39, 8'd136, 8'd85, 8'd97, 8'd103, 8'd108, 8'd184, 8'd192, 8'd196, 8'd194, 8'd91, 8'd112, 8'd125, 8'd150, 8'd114, 8'd118, 8'd118, 8'd104, 8'd148, 8'd147, 8'd137, 8'd225, 8'd154, 8'd112, 8'd164, 8'd63, 8'd59, 8'd55, 8'd64, 8'd88, 8'd70, 8'd97, 8'd115, 8'd74, 8'd220, 8'd144, 8'd119, 8'd129, 8'd106, 8'd148, 8'd123, 8'd89, 8'd94, 8'd100, 8'd141, 8'd166, 8'd147, 8'd195, 8'd208, 8'd177, 8'd206, 8'd111, 8'd140, 8'd151, 8'd81, 8'd113, 8'd52, 8'd68, 8'd68, 8'd82, 8'd110, 8'd141, 8'd164, 8'd174, 8'd89, 8'd77, 8'd131, 8'd119, 8'd90, 8'd95, 8'd120, 8'd98, 8'd92, 8'd150, 8'd153, 8'd146, 8'd230, 8'd138, 8'd207, 8'd131, 8'd105, 8'd136, 8'd115, 8'd41, 8'd137, 8'd136, 8'd80, 8'd154, 8'd163, 8'd111, 8'd213, 8'd137, 8'd161, 8'd123, 8'd79, 8'd74, 8'd86, 8'd93, 8'd105, 8'd68, 8'd157, 8'd128, 8'd161, 8'd145, 8'd225, 8'd149, 8'd168, 8'd188, 8'd160, 8'd136, 8'd117, 8'd99, 8'd58, 8'd56, 8'd132, 8'd124, 8'd174, 8'd141, 8'd127, 8'd169, 8'd95, 8'd90, 8'd145, 8'd71, 8'd71, 8'd50, 8'd49, 8'd160, 8'd147, 8'd138, 8'd105, 8'd164, 8'd139, 8'd214, 8'd167, 8'd153, 8'd144, 8'd162, 8'd97, 8'd83, 8'd85, 8'd70, 8'd92, 8'd105, 8'd175, 8'd130, 8'd170, 8'd164, 8'd117, 8'd119, 8'd92, 8'd137, 8'd99, 8'd89, 8'd56, 8'd128, 8'd79, 8'd126, 8'd158, 8'd137, 8'd220, 8'd150, 8'd124, 8'd155, 8'd157, 8'd140, 8'd158, 8'd49, 8'd142, 8'd128, 8'd101, 8'd90, 8'd93, 8'd152, 8'd155, 8'd131, 8'd140, 8'd116, 8'd163, 8'd139, 8'd75, 8'd132, 8'd135, 8'd94, 8'd116, 8'd72, 8'd114, 8'd169, 8'd129, 8'd131, 8'd118, 8'd151, 8'd114, 8'd127, 8'd127, 8'd132, 8'd83, 8'd58, 8'd115, 8'd96, 8'd136, 8'd102, 8'd93, 8'd147, 8'd161, 8'd120, 8'd126, 8'd70, 8'd50, 8'd29, 8'd102, 8'd116, 8'd41, 8'd68, 8'd86, 8'd166, 8'd134, 8'd93, 8'd96, 8'd64, 8'd91, 8'd99, 8'd133, 8'd46, 8'd68, 8'd41, 8'd70, 8'd148, 8'd151, 8'd36, 8'd90, 8'd132, 8'd121, 8'd125, 8'd132, 8'd48, 8'd39, 8'd85, 8'd50, 8'd40, 8'd69, 8'd100, 8'd86, 8'd126, 8'd104, 8'd166, 8'd71, 8'd133, 8'd141, 8'd74, 8'd134, 8'd48, 8'd102, 8'd49, 8'd111, 8'd135, 8'd101, 8'd67, 8'd97, 8'd65, 8'd148, 8'd147, 8'd71, 8'd87, 8'd39, 8'd110, 8'd38, 8'd89, 8'd98, 8'd115, 8'd142, 8'd115, 8'd108, 8'd156, 8'd161, 8'd127, 8'd93, 8'd124, 8'd50, 8'd129, 8'd97, 8'd89, 8'd94, 8'd89, 8'd59, 8'd131, 8'd42, 8'd110, 8'd123, 8'd83, 8'd103, 8'd91, 8'd81, 8'd97, 8'd41, 8'd91, 8'd97, 8'd88, 8'd88, 8'd135, 8'd60, 8'd77, 8'd138, 8'd79, 8'd106, 8'd70, 8'd129, 8'd125, 8'd90, 8'd144, 8'd99, 8'd67, 8'd90, 8'd128, 8'd119, 8'd109, 8'd117, 8'd114, 8'd100, 8'd62, 8'd61, 8'd95, 8'd50, 8'd130, 8'd89, 8'd69, 8'd108, 8'd77, 8'd77, 8'd137, 8'd103, 8'd70, 8'd99, 8'd108, 8'd74, 8'd102, 8'd112, 8'd133, 8'd71, 8'd98, 8'd134, 8'd57, 8'd105, 8'd107, 8'd132, 8'd111, 8'd117, 8'd114, 8'd65, 8'd90, 8'd104, 8'd67, 8'd121, 8'd89, 8'd135, 8'd67, 8'd48, 8'd88, 8'd85, 8'd114, 8'd87, 8'd110, 8'd90, 8'd96, 8'd44, 8'd155, 8'd64, 8'd101, 8'd133, 8'd148, 8'd143, 8'd126, 8'd113, 8'd139, 8'd142, 8'd79, 8'd165, 8'd150, 8'd105, 8'd84, 8'd134, 8'd108, 8'd99, 8'd109, 8'd85, 8'd70, 8'd69, 8'd122, 8'd126, 8'd98, 8'd121, 8'd112, 8'd45, 8'd114, 8'd96, 8'd122, 8'd77, 8'd157, 8'd85, 8'd142, 8'd166, 8'd112, 8'd150, 8'd178, 8'd191, 8'd187, 8'd110, 8'd160, 8'd137, 8'd94, 8'd111, 8'd93, 8'd112, 8'd114, 8'd129, 8'd161, 8'd106, 8'd61, 8'd73, 8'd135, 8'd67, 8'd161, 8'd78, 8'd119, 8'd83, 8'd84, 8'd107, 8'd137, 8'd127, 8'd129, 8'd180, 8'd164, 8'd156, 8'd156, 8'd209, 8'd184, 8'd126, 8'd174, 8'd110, 8'd163, 8'd108, 8'd125, 8'd114, 8'd89, 8'd110, 8'd151, 8'd144, 8'd132, 8'd127, 8'd139, 8'd104, 8'd101, 8'd136, 8'd80, 8'd123, 8'd124, 8'd118, 8'd197, 8'd168, 8'd187, 8'd158, 8'd172, 8'd180, 8'd186, 8'd132, 8'd107, 8'd153, 8'd136, 8'd139, 8'd167, 8'd213, 8'd106, 8'd148, 8'd142, 8'd153, 8'd154, 8'd119, 8'd103, 8'd160, 8'd150, 8'd149, 8'd139, 8'd109, 8'd104, 8'd170, 8'd201, 8'd166, 8'd175, 8'd198, 8'd181, 8'd158, 8'd182, 8'd142, 8'd124, 8'd143, 8'd189, 8'd166, 8'd142, 8'd146, 8'd177, 8'd184, 8'd170, 8'd128, 8'd128, 8'd172, 8'd78, 8'd165, 8'd77, 8'd124, 8'd121, 8'd125, 8'd115, 8'd120, 8'd144, 8'd125, 8'd153, 8'd146, 8'd167, 8'd147, 8'd186, 8'd163, 8'd160, 8'd189, 8'd107, 8'd127, 8'd150, 8'd98, 8'd91, 8'd119, 8'd98, 8'd87, 8'd137, 8'd141, 8'd97, 8'd98, 8'd115, 8'd106, 8'd149, 8'd88, 8'd115, 8'd133, 8'd133, 8'd118, 8'd123, 8'd71, 8'd151, 8'd152, 8'd74, 8'd70, 8'd166, 8'd87, 8'd176, 8'd162, 8'd160, 8'd141, 8'd115, 8'd139, 8'd81, 8'd149, 8'd75, 8'd122, 8'd84, 8'd113, 8'd123})
) cell_0_84 (
    .clk(clk),
    .input_index(index_0_83_84),
    .input_value(value_0_83_84),
    .input_result(result_0_83_84),
    .input_enable(enable_0_83_84),
    .output_index(index_0_84_85),
    .output_value(value_0_84_85),
    .output_result(result_0_84_85),
    .output_enable(enable_0_84_85)
);

wire [10-1:0] index_0_85_86;
wire [`DATA_WIDTH-1:0] value_0_85_86;
wire [`DATA_WIDTH*4:0] result_0_85_86;
wire enable_0_85_86;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd126, 8'd159, 8'd129, 8'd138, 8'd63, 8'd82, 8'd115, 8'd98, 8'd149, 8'd134, 8'd91, 8'd57, 8'd98, 8'd138, 8'd89, 8'd80, 8'd144, 8'd141, 8'd105, 8'd60, 8'd61, 8'd101, 8'd102, 8'd97, 8'd75, 8'd135, 8'd161, 8'd76, 8'd76, 8'd97, 8'd125, 8'd86, 8'd124, 8'd123, 8'd88, 8'd75, 8'd73, 8'd133, 8'd111, 8'd60, 8'd77, 8'd62, 8'd97, 8'd119, 8'd146, 8'd154, 8'd73, 8'd106, 8'd94, 8'd152, 8'd161, 8'd179, 8'd169, 8'd104, 8'd159, 8'd115, 8'd138, 8'd138, 8'd157, 8'd154, 8'd150, 8'd53, 8'd126, 8'd165, 8'd88, 8'd75, 8'd97, 8'd118, 8'd68, 8'd126, 8'd152, 8'd60, 8'd79, 8'd104, 8'd154, 8'd155, 8'd107, 8'd111, 8'd163, 8'd105, 8'd80, 8'd153, 8'd95, 8'd141, 8'd139, 8'd165, 8'd122, 8'd169, 8'd108, 8'd120, 8'd190, 8'd152, 8'd143, 8'd84, 8'd153, 8'd127, 8'd93, 8'd182, 8'd104, 8'd97, 8'd142, 8'd174, 8'd159, 8'd127, 8'd91, 8'd129, 8'd130, 8'd134, 8'd69, 8'd105, 8'd73, 8'd138, 8'd90, 8'd113, 8'd165, 8'd80, 8'd116, 8'd129, 8'd137, 8'd122, 8'd142, 8'd151, 8'd129, 8'd86, 8'd146, 8'd176, 8'd160, 8'd142, 8'd148, 8'd171, 8'd82, 8'd151, 8'd144, 8'd156, 8'd153, 8'd62, 8'd118, 8'd81, 8'd114, 8'd143, 8'd120, 8'd89, 8'd139, 8'd133, 8'd109, 8'd167, 8'd115, 8'd92, 8'd107, 8'd131, 8'd145, 8'd149, 8'd145, 8'd67, 8'd83, 8'd86, 8'd114, 8'd100, 8'd93, 8'd116, 8'd103, 8'd164, 8'd102, 8'd164, 8'd85, 8'd110, 8'd159, 8'd160, 8'd154, 8'd79, 8'd165, 8'd90, 8'd142, 8'd79, 8'd108, 8'd110, 8'd168, 8'd111, 8'd146, 8'd150, 8'd123, 8'd133, 8'd79, 8'd124, 8'd111, 8'd83, 8'd114, 8'd162, 8'd126, 8'd84, 8'd74, 8'd169, 8'd105, 8'd145, 8'd79, 8'd100, 8'd102, 8'd93, 8'd124, 8'd102, 8'd159, 8'd144, 8'd143, 8'd75, 8'd150, 8'd122, 8'd148, 8'd127, 8'd62, 8'd69, 8'd83, 8'd112, 8'd128, 8'd88, 8'd141, 8'd129, 8'd87, 8'd73, 8'd106, 8'd102, 8'd94, 8'd123, 8'd102, 8'd152, 8'd165, 8'd96, 8'd114, 8'd164, 8'd103, 8'd73, 8'd127, 8'd92, 8'd147, 8'd138, 8'd153, 8'd149, 8'd145, 8'd94, 8'd133, 8'd108, 8'd100, 8'd99, 8'd155, 8'd135, 8'd83, 8'd107, 8'd80, 8'd90, 8'd141, 8'd96, 8'd82, 8'd123, 8'd101, 8'd169, 8'd111, 8'd174, 8'd148, 8'd122, 8'd76, 8'd128, 8'd148, 8'd140, 8'd159, 8'd181, 8'd117, 8'd170, 8'd77, 8'd167, 8'd150, 8'd131, 8'd108, 8'd114, 8'd164, 8'd80, 8'd88, 8'd121, 8'd124, 8'd98, 8'd114, 8'd95, 8'd135, 8'd109, 8'd191, 8'd160, 8'd77, 8'd135, 8'd72, 8'd112, 8'd126, 8'd116, 8'd142, 8'd148, 8'd167, 8'd132, 8'd141, 8'd147, 8'd159, 8'd147, 8'd178, 8'd112, 8'd146, 8'd76, 8'd98, 8'd102, 8'd155, 8'd111, 8'd140, 8'd133, 8'd116, 8'd179, 8'd139, 8'd102, 8'd62, 8'd136, 8'd145, 8'd127, 8'd117, 8'd138, 8'd183, 8'd124, 8'd157, 8'd109, 8'd179, 8'd163, 8'd151, 8'd101, 8'd149, 8'd154, 8'd148, 8'd167, 8'd131, 8'd179, 8'd130, 8'd78, 8'd108, 8'd133, 8'd154, 8'd129, 8'd133, 8'd72, 8'd142, 8'd141, 8'd72, 8'd133, 8'd104, 8'd126, 8'd131, 8'd108, 8'd140, 8'd101, 8'd121, 8'd109, 8'd143, 8'd124, 8'd85, 8'd119, 8'd98, 8'd180, 8'd134, 8'd159, 8'd139, 8'd152, 8'd135, 8'd90, 8'd181, 8'd130, 8'd117, 8'd120, 8'd82, 8'd152, 8'd75, 8'd95, 8'd110, 8'd107, 8'd135, 8'd172, 8'd118, 8'd129, 8'd69, 8'd129, 8'd147, 8'd89, 8'd101, 8'd98, 8'd102, 8'd163, 8'd62, 8'd127, 8'd111, 8'd119, 8'd115, 8'd104, 8'd159, 8'd128, 8'd152, 8'd129, 8'd70, 8'd159, 8'd96, 8'd132, 8'd102, 8'd102, 8'd139, 8'd148, 8'd169, 8'd109, 8'd89, 8'd153, 8'd86, 8'd117, 8'd160, 8'd90, 8'd102, 8'd75, 8'd100, 8'd127, 8'd71, 8'd129, 8'd125, 8'd128, 8'd108, 8'd133, 8'd90, 8'd172, 8'd71, 8'd105, 8'd160, 8'd166, 8'd182, 8'd147, 8'd156, 8'd124, 8'd116, 8'd92, 8'd40, 8'd93, 8'd98, 8'd151, 8'd125, 8'd97, 8'd99, 8'd60, 8'd90, 8'd91, 8'd73, 8'd138, 8'd83, 8'd154, 8'd74, 8'd136, 8'd126, 8'd111, 8'd66, 8'd143, 8'd166, 8'd123, 8'd110, 8'd148, 8'd105, 8'd180, 8'd151, 8'd63, 8'd89, 8'd101, 8'd65, 8'd96, 8'd120, 8'd72, 8'd118, 8'd115, 8'd115, 8'd147, 8'd120, 8'd73, 8'd66, 8'd76, 8'd132, 8'd47, 8'd62, 8'd99, 8'd71, 8'd98, 8'd183, 8'd111, 8'd147, 8'd115, 8'd182, 8'd178, 8'd138, 8'd106, 8'd113, 8'd107, 8'd94, 8'd75, 8'd107, 8'd95, 8'd163, 8'd146, 8'd165, 8'd148, 8'd70, 8'd86, 8'd118, 8'd87, 8'd88, 8'd65, 8'd112, 8'd13, 8'd81, 8'd123, 8'd109, 8'd113, 8'd116, 8'd157, 8'd191, 8'd148, 8'd104, 8'd94, 8'd153, 8'd131, 8'd140, 8'd116, 8'd119, 8'd160, 8'd144, 8'd133, 8'd102, 8'd167, 8'd151, 8'd134, 8'd154, 8'd102, 8'd143, 8'd143, 8'd108, 8'd66, 8'd69, 8'd111, 8'd108, 8'd170, 8'd151, 8'd91, 8'd93, 8'd102, 8'd174, 8'd166, 8'd149, 8'd97, 8'd141, 8'd117, 8'd104, 8'd108, 8'd93, 8'd137, 8'd184, 8'd133, 8'd165, 8'd161, 8'd147, 8'd130, 8'd141, 8'd127, 8'd67, 8'd57, 8'd140, 8'd168, 8'd100, 8'd170, 8'd121, 8'd77, 8'd132, 8'd100, 8'd86, 8'd155, 8'd98, 8'd71, 8'd153, 8'd137, 8'd101, 8'd138, 8'd115, 8'd156, 8'd114, 8'd159, 8'd129, 8'd100, 8'd70, 8'd103, 8'd123, 8'd146, 8'd143, 8'd98, 8'd138, 8'd124, 8'd145, 8'd64, 8'd103, 8'd118, 8'd110, 8'd160, 8'd157, 8'd151, 8'd108, 8'd136, 8'd175, 8'd88, 8'd96, 8'd177, 8'd131, 8'd106, 8'd134, 8'd136, 8'd98, 8'd125, 8'd81, 8'd102, 8'd80, 8'd52, 8'd87, 8'd103, 8'd130, 8'd72, 8'd73, 8'd58, 8'd99, 8'd68, 8'd107, 8'd121, 8'd95, 8'd163, 8'd104, 8'd93, 8'd108, 8'd109, 8'd104, 8'd163, 8'd176, 8'd113, 8'd160, 8'd168, 8'd82, 8'd106, 8'd136, 8'd130, 8'd80, 8'd120, 8'd94, 8'd126, 8'd82, 8'd35, 8'd85, 8'd122, 8'd87, 8'd83, 8'd65, 8'd109, 8'd128, 8'd130, 8'd134, 8'd112, 8'd158, 8'd75, 8'd78, 8'd85, 8'd136, 8'd115, 8'd95, 8'd70, 8'd110, 8'd105, 8'd145, 8'd75, 8'd97, 8'd97, 8'd147, 8'd100, 8'd122, 8'd102, 8'd79, 8'd122, 8'd124, 8'd54, 8'd132, 8'd95, 8'd90, 8'd51, 8'd97, 8'd96, 8'd96, 8'd134, 8'd118, 8'd103, 8'd91, 8'd143, 8'd169, 8'd105, 8'd65, 8'd91, 8'd114, 8'd168, 8'd87, 8'd90, 8'd130, 8'd133, 8'd67, 8'd126, 8'd60, 8'd74, 8'd108, 8'd122, 8'd124, 8'd93, 8'd130, 8'd120, 8'd121, 8'd114, 8'd96, 8'd143, 8'd121, 8'd138, 8'd127, 8'd80, 8'd162, 8'd98, 8'd147, 8'd82, 8'd91, 8'd143, 8'd109, 8'd164, 8'd82, 8'd160, 8'd157, 8'd76, 8'd63, 8'd124, 8'd145, 8'd62, 8'd84, 8'd119, 8'd146, 8'd151, 8'd133, 8'd120, 8'd132, 8'd66, 8'd103, 8'd84, 8'd81, 8'd80, 8'd100, 8'd129, 8'd159, 8'd154, 8'd169, 8'd102, 8'd106, 8'd113, 8'd105, 8'd91, 8'd98, 8'd130, 8'd107, 8'd163, 8'd162, 8'd134, 8'd141, 8'd105, 8'd82, 8'd119, 8'd120, 8'd68, 8'd132, 8'd146, 8'd79, 8'd157, 8'd86, 8'd87, 8'd145, 8'd96, 8'd161, 8'd97, 8'd117, 8'd110})
) cell_0_85 (
    .clk(clk),
    .input_index(index_0_84_85),
    .input_value(value_0_84_85),
    .input_result(result_0_84_85),
    .input_enable(enable_0_84_85),
    .output_index(index_0_85_86),
    .output_value(value_0_85_86),
    .output_result(result_0_85_86),
    .output_enable(enable_0_85_86)
);

wire [10-1:0] index_0_86_87;
wire [`DATA_WIDTH-1:0] value_0_86_87;
wire [`DATA_WIDTH*4:0] result_0_86_87;
wire enable_0_86_87;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd103, 8'd131, 8'd113, 8'd99, 8'd144, 8'd128, 8'd162, 8'd139, 8'd102, 8'd183, 8'd195, 8'd92, 8'd148, 8'd140, 8'd164, 8'd140, 8'd116, 8'd142, 8'd91, 8'd185, 8'd175, 8'd147, 8'd163, 8'd130, 8'd116, 8'd89, 8'd114, 8'd160, 8'd115, 8'd86, 8'd151, 8'd120, 8'd74, 8'd132, 8'd136, 8'd128, 8'd129, 8'd98, 8'd97, 8'd77, 8'd115, 8'd113, 8'd93, 8'd67, 8'd85, 8'd100, 8'd121, 8'd140, 8'd145, 8'd146, 8'd68, 8'd62, 8'd114, 8'd117, 8'd160, 8'd96, 8'd95, 8'd81, 8'd85, 8'd61, 8'd100, 8'd131, 8'd123, 8'd132, 8'd73, 8'd78, 8'd121, 8'd94, 8'd86, 8'd132, 8'd108, 8'd90, 8'd136, 8'd142, 8'd114, 8'd150, 8'd135, 8'd72, 8'd127, 8'd152, 8'd135, 8'd139, 8'd89, 8'd164, 8'd117, 8'd117, 8'd132, 8'd94, 8'd28, 8'd80, 8'd52, 8'd58, 8'd120, 8'd122, 8'd152, 8'd148, 8'd138, 8'd108, 8'd133, 8'd177, 8'd79, 8'd108, 8'd143, 8'd112, 8'd80, 8'd123, 8'd97, 8'd131, 8'd149, 8'd128, 8'd152, 8'd78, 8'd93, 8'd84, 8'd56, 8'd53, 8'd71, 8'd111, 8'd143, 8'd74, 8'd75, 8'd161, 8'd160, 8'd90, 8'd166, 8'd131, 8'd83, 8'd159, 8'd76, 8'd139, 8'd112, 8'd138, 8'd156, 8'd132, 8'd143, 8'd76, 8'd152, 8'd82, 8'd121, 8'd97, 8'd92, 8'd82, 8'd97, 8'd89, 8'd67, 8'd142, 8'd65, 8'd151, 8'd161, 8'd110, 8'd86, 8'd143, 8'd162, 8'd88, 8'd158, 8'd91, 8'd74, 8'd108, 8'd156, 8'd82, 8'd80, 8'd122, 8'd106, 8'd138, 8'd78, 8'd169, 8'd146, 8'd141, 8'd165, 8'd141, 8'd127, 8'd62, 8'd104, 8'd84, 8'd104, 8'd165, 8'd125, 8'd155, 8'd77, 8'd154, 8'd110, 8'd142, 8'd91, 8'd139, 8'd92, 8'd135, 8'd122, 8'd131, 8'd85, 8'd147, 8'd164, 8'd148, 8'd97, 8'd149, 8'd80, 8'd140, 8'd120, 8'd164, 8'd118, 8'd134, 8'd151, 8'd126, 8'd147, 8'd152, 8'd77, 8'd92, 8'd117, 8'd137, 8'd124, 8'd148, 8'd124, 8'd106, 8'd98, 8'd124, 8'd163, 8'd109, 8'd83, 8'd124, 8'd105, 8'd139, 8'd78, 8'd70, 8'd130, 8'd134, 8'd158, 8'd100, 8'd85, 8'd84, 8'd70, 8'd152, 8'd108, 8'd119, 8'd171, 8'd79, 8'd122, 8'd154, 8'd116, 8'd97, 8'd124, 8'd104, 8'd138, 8'd172, 8'd91, 8'd145, 8'd145, 8'd149, 8'd93, 8'd130, 8'd102, 8'd147, 8'd123, 8'd168, 8'd142, 8'd116, 8'd61, 8'd85, 8'd98, 8'd162, 8'd77, 8'd78, 8'd162, 8'd176, 8'd114, 8'd73, 8'd113, 8'd74, 8'd111, 8'd101, 8'd119, 8'd126, 8'd93, 8'd87, 8'd148, 8'd82, 8'd70, 8'd83, 8'd158, 8'd97, 8'd108, 8'd93, 8'd92, 8'd145, 8'd69, 8'd153, 8'd177, 8'd163, 8'd81, 8'd157, 8'd135, 8'd134, 8'd142, 8'd154, 8'd150, 8'd117, 8'd163, 8'd176, 8'd184, 8'd163, 8'd103, 8'd103, 8'd119, 8'd95, 8'd116, 8'd106, 8'd125, 8'd125, 8'd174, 8'd129, 8'd150, 8'd92, 8'd153, 8'd124, 8'd132, 8'd139, 8'd96, 8'd137, 8'd97, 8'd160, 8'd150, 8'd115, 8'd109, 8'd143, 8'd104, 8'd131, 8'd91, 8'd96, 8'd113, 8'd132, 8'd83, 8'd96, 8'd162, 8'd137, 8'd116, 8'd156, 8'd170, 8'd146, 8'd73, 8'd125, 8'd120, 8'd140, 8'd114, 8'd98, 8'd144, 8'd75, 8'd90, 8'd109, 8'd140, 8'd98, 8'd173, 8'd152, 8'd146, 8'd87, 8'd124, 8'd93, 8'd115, 8'd118, 8'd160, 8'd111, 8'd102, 8'd88, 8'd150, 8'd94, 8'd114, 8'd113, 8'd160, 8'd55, 8'd101, 8'd130, 8'd133, 8'd136, 8'd93, 8'd64, 8'd107, 8'd68, 8'd88, 8'd161, 8'd89, 8'd138, 8'd107, 8'd131, 8'd123, 8'd94, 8'd150, 8'd141, 8'd98, 8'd158, 8'd160, 8'd96, 8'd155, 8'd177, 8'd118, 8'd71, 8'd142, 8'd131, 8'd110, 8'd119, 8'd212, 8'd183, 8'd160, 8'd103, 8'd83, 8'd75, 8'd125, 8'd101, 8'd143, 8'd103, 8'd80, 8'd79, 8'd136, 8'd154, 8'd162, 8'd121, 8'd120, 8'd82, 8'd68, 8'd122, 8'd179, 8'd121, 8'd90, 8'd135, 8'd104, 8'd111, 8'd168, 8'd161, 8'd133, 8'd158, 8'd156, 8'd85, 8'd97, 8'd81, 8'd96, 8'd87, 8'd109, 8'd130, 8'd169, 8'd87, 8'd135, 8'd116, 8'd85, 8'd149, 8'd174, 8'd85, 8'd79, 8'd126, 8'd96, 8'd182, 8'd152, 8'd82, 8'd94, 8'd67, 8'd116, 8'd95, 8'd148, 8'd143, 8'd105, 8'd117, 8'd109, 8'd130, 8'd137, 8'd127, 8'd164, 8'd165, 8'd112, 8'd90, 8'd167, 8'd90, 8'd172, 8'd129, 8'd109, 8'd136, 8'd134, 8'd123, 8'd158, 8'd187, 8'd170, 8'd113, 8'd125, 8'd99, 8'd83, 8'd59, 8'd139, 8'd157, 8'd143, 8'd144, 8'd124, 8'd94, 8'd115, 8'd113, 8'd143, 8'd82, 8'd157, 8'd80, 8'd117, 8'd107, 8'd77, 8'd91, 8'd143, 8'd157, 8'd163, 8'd162, 8'd193, 8'd117, 8'd181, 8'd154, 8'd106, 8'd146, 8'd79, 8'd47, 8'd163, 8'd135, 8'd105, 8'd166, 8'd154, 8'd153, 8'd95, 8'd123, 8'd169, 8'd149, 8'd127, 8'd150, 8'd99, 8'd74, 8'd138, 8'd112, 8'd154, 8'd176, 8'd91, 8'd155, 8'd128, 8'd144, 8'd173, 8'd149, 8'd92, 8'd120, 8'd82, 8'd125, 8'd80, 8'd96, 8'd123, 8'd80, 8'd73, 8'd89, 8'd97, 8'd156, 8'd74, 8'd134, 8'd129, 8'd165, 8'd148, 8'd70, 8'd161, 8'd161, 8'd179, 8'd167, 8'd102, 8'd142, 8'd179, 8'd112, 8'd139, 8'd84, 8'd73, 8'd115, 8'd105, 8'd100, 8'd167, 8'd132, 8'd149, 8'd117, 8'd98, 8'd71, 8'd67, 8'd131, 8'd94, 8'd84, 8'd80, 8'd121, 8'd129, 8'd158, 8'd165, 8'd105, 8'd93, 8'd92, 8'd90, 8'd160, 8'd177, 8'd135, 8'd138, 8'd109, 8'd144, 8'd149, 8'd115, 8'd101, 8'd150, 8'd131, 8'd117, 8'd170, 8'd154, 8'd115, 8'd88, 8'd144, 8'd121, 8'd143, 8'd69, 8'd111, 8'd127, 8'd118, 8'd130, 8'd87, 8'd179, 8'd161, 8'd95, 8'd113, 8'd126, 8'd75, 8'd124, 8'd79, 8'd92, 8'd115, 8'd139, 8'd87, 8'd104, 8'd102, 8'd110, 8'd140, 8'd138, 8'd118, 8'd133, 8'd159, 8'd139, 8'd98, 8'd117, 8'd103, 8'd121, 8'd91, 8'd113, 8'd163, 8'd154, 8'd145, 8'd85, 8'd95, 8'd123, 8'd149, 8'd93, 8'd154, 8'd147, 8'd122, 8'd114, 8'd78, 8'd151, 8'd87, 8'd113, 8'd153, 8'd98, 8'd82, 8'd94, 8'd151, 8'd138, 8'd148, 8'd163, 8'd88, 8'd97, 8'd91, 8'd115, 8'd159, 8'd167, 8'd143, 8'd107, 8'd118, 8'd135, 8'd172, 8'd149, 8'd103, 8'd126, 8'd106, 8'd89, 8'd163, 8'd167, 8'd144, 8'd172, 8'd122, 8'd95, 8'd176, 8'd94, 8'd162, 8'd129, 8'd176, 8'd160, 8'd118, 8'd162, 8'd117, 8'd111, 8'd168, 8'd188, 8'd139, 8'd177, 8'd141, 8'd160, 8'd125, 8'd154, 8'd157, 8'd158, 8'd78, 8'd166, 8'd78, 8'd91, 8'd135, 8'd153, 8'd161, 8'd152, 8'd154, 8'd109, 8'd160, 8'd157, 8'd122, 8'd177, 8'd174, 8'd112, 8'd151, 8'd181, 8'd158, 8'd151, 8'd121, 8'd119, 8'd122, 8'd97, 8'd114, 8'd100, 8'd133, 8'd95, 8'd168, 8'd134, 8'd127, 8'd120, 8'd146, 8'd133, 8'd162, 8'd149, 8'd176, 8'd105, 8'd177, 8'd101, 8'd161, 8'd153, 8'd114, 8'd155, 8'd172, 8'd174, 8'd104, 8'd142, 8'd177, 8'd145, 8'd104, 8'd117, 8'd104, 8'd162, 8'd126, 8'd83, 8'd126, 8'd116, 8'd133, 8'd135, 8'd75, 8'd118, 8'd117, 8'd139, 8'd84, 8'd116, 8'd125, 8'd107, 8'd103, 8'd111, 8'd137, 8'd106, 8'd142, 8'd156, 8'd132, 8'd94, 8'd73, 8'd148, 8'd85, 8'd120, 8'd138, 8'd169, 8'd164})
) cell_0_86 (
    .clk(clk),
    .input_index(index_0_85_86),
    .input_value(value_0_85_86),
    .input_result(result_0_85_86),
    .input_enable(enable_0_85_86),
    .output_index(index_0_86_87),
    .output_value(value_0_86_87),
    .output_result(result_0_86_87),
    .output_enable(enable_0_86_87)
);

wire [10-1:0] index_0_87_88;
wire [`DATA_WIDTH-1:0] value_0_87_88;
wire [`DATA_WIDTH*4:0] result_0_87_88;
wire enable_0_87_88;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd141, 8'd102, 8'd127, 8'd98, 8'd156, 8'd165, 8'd117, 8'd184, 8'd104, 8'd96, 8'd183, 8'd102, 8'd121, 8'd147, 8'd101, 8'd160, 8'd178, 8'd154, 8'd96, 8'd146, 8'd149, 8'd123, 8'd105, 8'd98, 8'd165, 8'd76, 8'd156, 8'd111, 8'd80, 8'd98, 8'd133, 8'd162, 8'd117, 8'd143, 8'd146, 8'd180, 8'd159, 8'd181, 8'd191, 8'd181, 8'd176, 8'd224, 8'd160, 8'd133, 8'd164, 8'd144, 8'd178, 8'd193, 8'd187, 8'd179, 8'd164, 8'd178, 8'd151, 8'd104, 8'd83, 8'd155, 8'd119, 8'd84, 8'd148, 8'd173, 8'd152, 8'd140, 8'd151, 8'd166, 8'd164, 8'd160, 8'd168, 8'd128, 8'd176, 8'd176, 8'd166, 8'd135, 8'd190, 8'd197, 8'd202, 8'd147, 8'd197, 8'd204, 8'd133, 8'd150, 8'd181, 8'd114, 8'd118, 8'd140, 8'd136, 8'd142, 8'd76, 8'd98, 8'd91, 8'd112, 8'd74, 8'd126, 8'd130, 8'd56, 8'd79, 8'd134, 8'd79, 8'd120, 8'd85, 8'd98, 8'd73, 8'd120, 8'd88, 8'd150, 8'd175, 8'd120, 8'd173, 8'd158, 8'd131, 8'd127, 8'd139, 8'd70, 8'd125, 8'd168, 8'd144, 8'd150, 8'd136, 8'd135, 8'd141, 8'd122, 8'd72, 8'd43, 8'd139, 8'd116, 8'd106, 8'd123, 8'd115, 8'd150, 8'd61, 8'd104, 8'd111, 8'd95, 8'd119, 8'd145, 8'd109, 8'd117, 8'd82, 8'd107, 8'd104, 8'd119, 8'd129, 8'd89, 8'd117, 8'd106, 8'd139, 8'd71, 8'd108, 8'd86, 8'd57, 8'd112, 8'd97, 8'd129, 8'd92, 8'd76, 8'd125, 8'd135, 8'd144, 8'd81, 8'd132, 8'd73, 8'd116, 8'd147, 8'd79, 8'd85, 8'd127, 8'd126, 8'd73, 8'd139, 8'd105, 8'd86, 8'd98, 8'd63, 8'd113, 8'd80, 8'd132, 8'd117, 8'd52, 8'd109, 8'd134, 8'd148, 8'd174, 8'd110, 8'd157, 8'd155, 8'd106, 8'd79, 8'd59, 8'd129, 8'd152, 8'd60, 8'd117, 8'd136, 8'd57, 8'd108, 8'd77, 8'd125, 8'd169, 8'd149, 8'd137, 8'd143, 8'd98, 8'd83, 8'd63, 8'd149, 8'd141, 8'd143, 8'd166, 8'd138, 8'd164, 8'd159, 8'd151, 8'd116, 8'd159, 8'd139, 8'd150, 8'd141, 8'd115, 8'd121, 8'd161, 8'd100, 8'd111, 8'd113, 8'd114, 8'd88, 8'd83, 8'd133, 8'd57, 8'd126, 8'd130, 8'd123, 8'd63, 8'd146, 8'd106, 8'd134, 8'd78, 8'd141, 8'd143, 8'd106, 8'd100, 8'd113, 8'd146, 8'd109, 8'd151, 8'd94, 8'd126, 8'd101, 8'd75, 8'd118, 8'd128, 8'd165, 8'd101, 8'd149, 8'd92, 8'd86, 8'd107, 8'd77, 8'd72, 8'd124, 8'd161, 8'd137, 8'd172, 8'd124, 8'd81, 8'd138, 8'd67, 8'd65, 8'd69, 8'd94, 8'd89, 8'd99, 8'd145, 8'd102, 8'd74, 8'd139, 8'd131, 8'd81, 8'd100, 8'd80, 8'd154, 8'd141, 8'd95, 8'd111, 8'd112, 8'd111, 8'd144, 8'd131, 8'd80, 8'd144, 8'd116, 8'd145, 8'd162, 8'd59, 8'd104, 8'd72, 8'd116, 8'd104, 8'd160, 8'd116, 8'd117, 8'd95, 8'd128, 8'd102, 8'd163, 8'd98, 8'd78, 8'd68, 8'd169, 8'd104, 8'd153, 8'd83, 8'd121, 8'd85, 8'd76, 8'd135, 8'd123, 8'd167, 8'd125, 8'd105, 8'd124, 8'd140, 8'd63, 8'd66, 8'd104, 8'd128, 8'd160, 8'd125, 8'd131, 8'd169, 8'd181, 8'd173, 8'd98, 8'd151, 8'd65, 8'd153, 8'd140, 8'd102, 8'd144, 8'd31, 8'd106, 8'd76, 8'd91, 8'd186, 8'd168, 8'd176, 8'd157, 8'd123, 8'd114, 8'd82, 8'd46, 8'd33, 8'd60, 8'd56, 8'd86, 8'd133, 8'd162, 8'd130, 8'd176, 8'd136, 8'd92, 8'd143, 8'd62, 8'd87, 8'd77, 8'd82, 8'd83, 8'd67, 8'd88, 8'd138, 8'd102, 8'd122, 8'd99, 8'd145, 8'd149, 8'd142, 8'd150, 8'd113, 8'd130, 8'd85, 8'd88, 8'd114, 8'd169, 8'd125, 8'd111, 8'd137, 8'd155, 8'd192, 8'd186, 8'd133, 8'd79, 8'd175, 8'd104, 8'd129, 8'd141, 8'd107, 8'd104, 8'd165, 8'd120, 8'd162, 8'd113, 8'd121, 8'd145, 8'd82, 8'd104, 8'd93, 8'd128, 8'd97, 8'd42, 8'd83, 8'd88, 8'd121, 8'd143, 8'd128, 8'd156, 8'd119, 8'd162, 8'd123, 8'd142, 8'd148, 8'd148, 8'd99, 8'd104, 8'd131, 8'd132, 8'd167, 8'd165, 8'd96, 8'd166, 8'd109, 8'd85, 8'd151, 8'd163, 8'd132, 8'd94, 8'd100, 8'd129, 8'd166, 8'd128, 8'd102, 8'd111, 8'd158, 8'd124, 8'd106, 8'd96, 8'd148, 8'd129, 8'd160, 8'd125, 8'd121, 8'd95, 8'd48, 8'd74, 8'd72, 8'd110, 8'd166, 8'd130, 8'd175, 8'd75, 8'd152, 8'd96, 8'd126, 8'd55, 8'd90, 8'd131, 8'd101, 8'd152, 8'd118, 8'd167, 8'd75, 8'd86, 8'd96, 8'd127, 8'd142, 8'd137, 8'd114, 8'd140, 8'd91, 8'd151, 8'd71, 8'd52, 8'd104, 8'd151, 8'd97, 8'd66, 8'd107, 8'd77, 8'd90, 8'd69, 8'd86, 8'd122, 8'd115, 8'd92, 8'd152, 8'd85, 8'd142, 8'd148, 8'd122, 8'd91, 8'd60, 8'd116, 8'd86, 8'd75, 8'd93, 8'd89, 8'd165, 8'd95, 8'd72, 8'd117, 8'd82, 8'd105, 8'd119, 8'd54, 8'd146, 8'd66, 8'd93, 8'd134, 8'd141, 8'd130, 8'd105, 8'd85, 8'd101, 8'd80, 8'd60, 8'd91, 8'd54, 8'd77, 8'd71, 8'd140, 8'd107, 8'd135, 8'd99, 8'd141, 8'd165, 8'd117, 8'd75, 8'd30, 8'd93, 8'd135, 8'd66, 8'd83, 8'd119, 8'd141, 8'd95, 8'd94, 8'd113, 8'd196, 8'd186, 8'd97, 8'd108, 8'd158, 8'd79, 8'd92, 8'd126, 8'd143, 8'd80, 8'd66, 8'd94, 8'd69, 8'd78, 8'd148, 8'd87, 8'd72, 8'd83, 8'd29, 8'd113, 8'd150, 8'd145, 8'd70, 8'd77, 8'd100, 8'd92, 8'd126, 8'd180, 8'd181, 8'd188, 8'd160, 8'd89, 8'd131, 8'd141, 8'd146, 8'd79, 8'd90, 8'd100, 8'd72, 8'd71, 8'd152, 8'd103, 8'd75, 8'd117, 8'd136, 8'd54, 8'd78, 8'd117, 8'd93, 8'd67, 8'd136, 8'd88, 8'd82, 8'd134, 8'd152, 8'd99, 8'd124, 8'd88, 8'd148, 8'd168, 8'd132, 8'd146, 8'd89, 8'd71, 8'd108, 8'd66, 8'd127, 8'd112, 8'd76, 8'd137, 8'd87, 8'd89, 8'd157, 8'd122, 8'd91, 8'd121, 8'd123, 8'd110, 8'd104, 8'd96, 8'd132, 8'd78, 8'd121, 8'd45, 8'd128, 8'd52, 8'd135, 8'd60, 8'd147, 8'd116, 8'd148, 8'd150, 8'd144, 8'd94, 8'd64, 8'd127, 8'd57, 8'd115, 8'd144, 8'd89, 8'd119, 8'd97, 8'd141, 8'd129, 8'd115, 8'd186, 8'd131, 8'd105, 8'd121, 8'd93, 8'd76, 8'd84, 8'd76, 8'd66, 8'd101, 8'd54, 8'd57, 8'd118, 8'd136, 8'd157, 8'd69, 8'd127, 8'd151, 8'd79, 8'd95, 8'd111, 8'd76, 8'd109, 8'd113, 8'd142, 8'd160, 8'd162, 8'd160, 8'd166, 8'd166, 8'd190, 8'd125, 8'd171, 8'd128, 8'd118, 8'd99, 8'd175, 8'd130, 8'd95, 8'd167, 8'd115, 8'd88, 8'd142, 8'd85, 8'd164, 8'd78, 8'd80, 8'd99, 8'd116, 8'd162, 8'd127, 8'd129, 8'd167, 8'd162, 8'd95, 8'd150, 8'd153, 8'd139, 8'd113, 8'd107, 8'd125, 8'd126, 8'd166, 8'd108, 8'd96, 8'd126, 8'd93, 8'd115, 8'd141, 8'd173, 8'd165, 8'd107, 8'd119, 8'd88, 8'd160, 8'd89, 8'd78, 8'd150, 8'd144, 8'd108, 8'd135, 8'd82, 8'd164, 8'd88, 8'd134, 8'd103, 8'd113, 8'd130, 8'd159, 8'd156, 8'd113, 8'd77, 8'd107, 8'd175, 8'd174, 8'd132, 8'd142, 8'd163, 8'd151, 8'd161, 8'd180, 8'd114, 8'd105, 8'd128, 8'd160, 8'd127, 8'd85, 8'd148, 8'd132, 8'd137, 8'd160, 8'd122, 8'd90, 8'd146, 8'd83, 8'd162, 8'd127, 8'd80, 8'd150, 8'd108, 8'd76, 8'd124, 8'd135, 8'd71, 8'd145, 8'd110, 8'd149, 8'd134, 8'd109, 8'd72, 8'd126, 8'd163, 8'd168, 8'd99, 8'd113})
) cell_0_87 (
    .clk(clk),
    .input_index(index_0_86_87),
    .input_value(value_0_86_87),
    .input_result(result_0_86_87),
    .input_enable(enable_0_86_87),
    .output_index(index_0_87_88),
    .output_value(value_0_87_88),
    .output_result(result_0_87_88),
    .output_enable(enable_0_87_88)
);

wire [10-1:0] index_0_88_89;
wire [`DATA_WIDTH-1:0] value_0_88_89;
wire [`DATA_WIDTH*4:0] result_0_88_89;
wire enable_0_88_89;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd109, 8'd76, 8'd107, 8'd163, 8'd150, 8'd73, 8'd148, 8'd92, 8'd112, 8'd119, 8'd61, 8'd69, 8'd140, 8'd95, 8'd93, 8'd106, 8'd135, 8'd139, 8'd84, 8'd139, 8'd127, 8'd161, 8'd80, 8'd154, 8'd153, 8'd72, 8'd96, 8'd84, 8'd145, 8'd142, 8'd101, 8'd117, 8'd96, 8'd120, 8'd139, 8'd90, 8'd130, 8'd73, 8'd96, 8'd165, 8'd68, 8'd116, 8'd132, 8'd169, 8'd155, 8'd122, 8'd82, 8'd128, 8'd144, 8'd123, 8'd145, 8'd111, 8'd140, 8'd110, 8'd165, 8'd80, 8'd106, 8'd109, 8'd120, 8'd117, 8'd164, 8'd114, 8'd94, 8'd116, 8'd173, 8'd171, 8'd87, 8'd78, 8'd111, 8'd154, 8'd156, 8'd160, 8'd69, 8'd125, 8'd145, 8'd156, 8'd162, 8'd125, 8'd144, 8'd149, 8'd103, 8'd165, 8'd87, 8'd131, 8'd110, 8'd164, 8'd152, 8'd178, 8'd150, 8'd170, 8'd181, 8'd158, 8'd144, 8'd116, 8'd153, 8'd98, 8'd106, 8'd85, 8'd135, 8'd83, 8'd128, 8'd67, 8'd92, 8'd79, 8'd83, 8'd83, 8'd76, 8'd83, 8'd123, 8'd118, 8'd129, 8'd169, 8'd132, 8'd115, 8'd92, 8'd166, 8'd169, 8'd191, 8'd190, 8'd97, 8'd181, 8'd91, 8'd158, 8'd94, 8'd74, 8'd99, 8'd99, 8'd67, 8'd123, 8'd53, 8'd59, 8'd88, 8'd88, 8'd145, 8'd117, 8'd108, 8'd68, 8'd158, 8'd138, 8'd98, 8'd98, 8'd136, 8'd177, 8'd177, 8'd124, 8'd127, 8'd160, 8'd173, 8'd91, 8'd145, 8'd163, 8'd89, 8'd77, 8'd143, 8'd118, 8'd59, 8'd106, 8'd78, 8'd161, 8'd88, 8'd107, 8'd147, 8'd159, 8'd96, 8'd104, 8'd104, 8'd150, 8'd87, 8'd129, 8'd90, 8'd91, 8'd144, 8'd128, 8'd178, 8'd94, 8'd107, 8'd142, 8'd145, 8'd138, 8'd102, 8'd159, 8'd65, 8'd149, 8'd68, 8'd135, 8'd143, 8'd168, 8'd92, 8'd135, 8'd158, 8'd109, 8'd105, 8'd151, 8'd77, 8'd114, 8'd137, 8'd114, 8'd113, 8'd122, 8'd165, 8'd177, 8'd97, 8'd93, 8'd170, 8'd160, 8'd176, 8'd122, 8'd135, 8'd69, 8'd144, 8'd102, 8'd67, 8'd72, 8'd153, 8'd132, 8'd134, 8'd92, 8'd167, 8'd146, 8'd81, 8'd112, 8'd113, 8'd103, 8'd123, 8'd161, 8'd87, 8'd167, 8'd172, 8'd184, 8'd155, 8'd88, 8'd89, 8'd160, 8'd91, 8'd142, 8'd140, 8'd90, 8'd79, 8'd133, 8'd110, 8'd84, 8'd137, 8'd72, 8'd151, 8'd138, 8'd88, 8'd151, 8'd112, 8'd115, 8'd138, 8'd109, 8'd150, 8'd131, 8'd173, 8'd140, 8'd130, 8'd127, 8'd132, 8'd153, 8'd90, 8'd147, 8'd112, 8'd128, 8'd71, 8'd81, 8'd152, 8'd117, 8'd126, 8'd159, 8'd89, 8'd97, 8'd120, 8'd166, 8'd120, 8'd112, 8'd98, 8'd71, 8'd69, 8'd107, 8'd135, 8'd97, 8'd151, 8'd156, 8'd99, 8'd154, 8'd78, 8'd118, 8'd78, 8'd110, 8'd143, 8'd126, 8'd121, 8'd80, 8'd136, 8'd173, 8'd153, 8'd96, 8'd105, 8'd73, 8'd103, 8'd89, 8'd129, 8'd80, 8'd97, 8'd88, 8'd115, 8'd152, 8'd132, 8'd159, 8'd112, 8'd143, 8'd136, 8'd139, 8'd128, 8'd136, 8'd151, 8'd137, 8'd109, 8'd128, 8'd99, 8'd149, 8'd138, 8'd147, 8'd157, 8'd123, 8'd135, 8'd113, 8'd114, 8'd76, 8'd136, 8'd99, 8'd88, 8'd135, 8'd121, 8'd135, 8'd133, 8'd84, 8'd106, 8'd98, 8'd84, 8'd139, 8'd87, 8'd99, 8'd109, 8'd131, 8'd134, 8'd107, 8'd142, 8'd155, 8'd174, 8'd193, 8'd161, 8'd107, 8'd151, 8'd81, 8'd139, 8'd124, 8'd122, 8'd74, 8'd126, 8'd162, 8'd107, 8'd75, 8'd129, 8'd135, 8'd83, 8'd150, 8'd56, 8'd112, 8'd91, 8'd82, 8'd128, 8'd61, 8'd66, 8'd105, 8'd170, 8'd152, 8'd207, 8'd122, 8'd194, 8'd147, 8'd147, 8'd145, 8'd97, 8'd97, 8'd160, 8'd131, 8'd81, 8'd85, 8'd93, 8'd135, 8'd130, 8'd109, 8'd122, 8'd103, 8'd94, 8'd112, 8'd96, 8'd143, 8'd109, 8'd161, 8'd103, 8'd168, 8'd107, 8'd195, 8'd167, 8'd221, 8'd145, 8'd106, 8'd106, 8'd129, 8'd110, 8'd113, 8'd76, 8'd131, 8'd114, 8'd113, 8'd127, 8'd127, 8'd84, 8'd105, 8'd142, 8'd105, 8'd55, 8'd52, 8'd90, 8'd139, 8'd110, 8'd119, 8'd149, 8'd153, 8'd89, 8'd142, 8'd206, 8'd204, 8'd124, 8'd77, 8'd95, 8'd97, 8'd148, 8'd129, 8'd124, 8'd139, 8'd105, 8'd92, 8'd69, 8'd97, 8'd99, 8'd145, 8'd127, 8'd156, 8'd94, 8'd139, 8'd98, 8'd107, 8'd76, 8'd107, 8'd115, 8'd141, 8'd71, 8'd161, 8'd166, 8'd109, 8'd88, 8'd156, 8'd73, 8'd162, 8'd108, 8'd127, 8'd116, 8'd144, 8'd76, 8'd139, 8'd102, 8'd70, 8'd123, 8'd59, 8'd165, 8'd149, 8'd129, 8'd102, 8'd61, 8'd74, 8'd119, 8'd49, 8'd93, 8'd122, 8'd117, 8'd140, 8'd118, 8'd158, 8'd117, 8'd118, 8'd151, 8'd70, 8'd92, 8'd97, 8'd139, 8'd75, 8'd60, 8'd60, 8'd41, 8'd151, 8'd102, 8'd147, 8'd166, 8'd107, 8'd52, 8'd32, 8'd48, 8'd105, 8'd112, 8'd44, 8'd76, 8'd75, 8'd132, 8'd114, 8'd83, 8'd129, 8'd163, 8'd96, 8'd118, 8'd60, 8'd78, 8'd67, 8'd132, 8'd86, 8'd118, 8'd42, 8'd91, 8'd86, 8'd143, 8'd93, 8'd108, 8'd124, 8'd146, 8'd102, 8'd66, 8'd139, 8'd54, 8'd47, 8'd57, 8'd63, 8'd150, 8'd83, 8'd99, 8'd163, 8'd154, 8'd129, 8'd122, 8'd117, 8'd55, 8'd64, 8'd125, 8'd34, 8'd114, 8'd69, 8'd89, 8'd119, 8'd149, 8'd108, 8'd127, 8'd166, 8'd154, 8'd53, 8'd125, 8'd91, 8'd71, 8'd83, 8'd89, 8'd150, 8'd96, 8'd175, 8'd144, 8'd139, 8'd103, 8'd119, 8'd111, 8'd100, 8'd116, 8'd87, 8'd107, 8'd59, 8'd79, 8'd115, 8'd59, 8'd76, 8'd144, 8'd95, 8'd129, 8'd142, 8'd92, 8'd64, 8'd112, 8'd57, 8'd154, 8'd141, 8'd129, 8'd121, 8'd78, 8'd91, 8'd86, 8'd98, 8'd106, 8'd85, 8'd105, 8'd76, 8'd49, 8'd76, 8'd66, 8'd90, 8'd81, 8'd47, 8'd135, 8'd67, 8'd121, 8'd119, 8'd182, 8'd184, 8'd98, 8'd104, 8'd137, 8'd120, 8'd154, 8'd123, 8'd143, 8'd121, 8'd126, 8'd109, 8'd111, 8'd146, 8'd182, 8'd87, 8'd86, 8'd54, 8'd123, 8'd138, 8'd100, 8'd138, 8'd122, 8'd96, 8'd104, 8'd128, 8'd115, 8'd143, 8'd155, 8'd142, 8'd163, 8'd101, 8'd139, 8'd125, 8'd105, 8'd105, 8'd148, 8'd156, 8'd164, 8'd144, 8'd164, 8'd140, 8'd128, 8'd144, 8'd136, 8'd151, 8'd149, 8'd124, 8'd105, 8'd134, 8'd140, 8'd85, 8'd154, 8'd144, 8'd146, 8'd138, 8'd110, 8'd168, 8'd156, 8'd163, 8'd179, 8'd169, 8'd173, 8'd90, 8'd156, 8'd78, 8'd132, 8'd158, 8'd130, 8'd73, 8'd121, 8'd120, 8'd150, 8'd146, 8'd82, 8'd109, 8'd97, 8'd134, 8'd104, 8'd127, 8'd117, 8'd112, 8'd109, 8'd139, 8'd94, 8'd130, 8'd70, 8'd87, 8'd93, 8'd72, 8'd127, 8'd153, 8'd163, 8'd114, 8'd106, 8'd168, 8'd168, 8'd92, 8'd135, 8'd75, 8'd101, 8'd155, 8'd97, 8'd123, 8'd157, 8'd77, 8'd139, 8'd152, 8'd94, 8'd166, 8'd107, 8'd118, 8'd147, 8'd121, 8'd138, 8'd78, 8'd86, 8'd109, 8'd149, 8'd128, 8'd135, 8'd101, 8'd142, 8'd95, 8'd106, 8'd129, 8'd63, 8'd153, 8'd131, 8'd75, 8'd159, 8'd112, 8'd155, 8'd160, 8'd139, 8'd83, 8'd132, 8'd82, 8'd115, 8'd83, 8'd76, 8'd91, 8'd149, 8'd112, 8'd71, 8'd115, 8'd104, 8'd72, 8'd132, 8'd129, 8'd148, 8'd123, 8'd97, 8'd76, 8'd112, 8'd160, 8'd80, 8'd136, 8'd164, 8'd134, 8'd124, 8'd124, 8'd155, 8'd71, 8'd86, 8'd149, 8'd78})
) cell_0_88 (
    .clk(clk),
    .input_index(index_0_87_88),
    .input_value(value_0_87_88),
    .input_result(result_0_87_88),
    .input_enable(enable_0_87_88),
    .output_index(index_0_88_89),
    .output_value(value_0_88_89),
    .output_result(result_0_88_89),
    .output_enable(enable_0_88_89)
);

wire [10-1:0] index_0_89_90;
wire [`DATA_WIDTH-1:0] value_0_89_90;
wire [`DATA_WIDTH*4:0] result_0_89_90;
wire enable_0_89_90;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd95, 8'd71, 8'd152, 8'd123, 8'd144, 8'd125, 8'd149, 8'd146, 8'd160, 8'd175, 8'd154, 8'd180, 8'd164, 8'd135, 8'd111, 8'd162, 8'd139, 8'd186, 8'd104, 8'd172, 8'd186, 8'd158, 8'd111, 8'd119, 8'd115, 8'd99, 8'd131, 8'd164, 8'd100, 8'd120, 8'd123, 8'd165, 8'd110, 8'd97, 8'd159, 8'd145, 8'd192, 8'd111, 8'd128, 8'd181, 8'd177, 8'd209, 8'd171, 8'd126, 8'd168, 8'd132, 8'd166, 8'd153, 8'd147, 8'd112, 8'd118, 8'd162, 8'd130, 8'd163, 8'd165, 8'd146, 8'd101, 8'd147, 8'd100, 8'd104, 8'd160, 8'd119, 8'd132, 8'd105, 8'd115, 8'd208, 8'd213, 8'd161, 8'd186, 8'd176, 8'd189, 8'd179, 8'd214, 8'd223, 8'd162, 8'd167, 8'd175, 8'd152, 8'd195, 8'd128, 8'd153, 8'd91, 8'd147, 8'd124, 8'd124, 8'd115, 8'd65, 8'd85, 8'd98, 8'd117, 8'd79, 8'd170, 8'd107, 8'd97, 8'd185, 8'd109, 8'd192, 8'd195, 8'd155, 8'd122, 8'd144, 8'd142, 8'd132, 8'd188, 8'd185, 8'd157, 8'd127, 8'd124, 8'd189, 8'd100, 8'd156, 8'd101, 8'd105, 8'd156, 8'd80, 8'd89, 8'd159, 8'd88, 8'd149, 8'd146, 8'd109, 8'd76, 8'd122, 8'd136, 8'd131, 8'd130, 8'd81, 8'd146, 8'd132, 8'd98, 8'd144, 8'd117, 8'd156, 8'd150, 8'd135, 8'd148, 8'd168, 8'd120, 8'd138, 8'd86, 8'd103, 8'd162, 8'd106, 8'd162, 8'd172, 8'd154, 8'd108, 8'd73, 8'd168, 8'd161, 8'd123, 8'd95, 8'd117, 8'd152, 8'd159, 8'd73, 8'd164, 8'd81, 8'd128, 8'd76, 8'd112, 8'd105, 8'd84, 8'd155, 8'd130, 8'd152, 8'd106, 8'd84, 8'd80, 8'd137, 8'd77, 8'd94, 8'd76, 8'd126, 8'd88, 8'd167, 8'd134, 8'd136, 8'd143, 8'd126, 8'd82, 8'd99, 8'd140, 8'd98, 8'd60, 8'd98, 8'd70, 8'd107, 8'd154, 8'd153, 8'd117, 8'd113, 8'd149, 8'd106, 8'd112, 8'd120, 8'd72, 8'd83, 8'd95, 8'd159, 8'd124, 8'd93, 8'd74, 8'd95, 8'd130, 8'd146, 8'd157, 8'd72, 8'd90, 8'd146, 8'd136, 8'd104, 8'd62, 8'd61, 8'd163, 8'd97, 8'd166, 8'd131, 8'd91, 8'd92, 8'd139, 8'd115, 8'd130, 8'd165, 8'd142, 8'd68, 8'd125, 8'd138, 8'd148, 8'd163, 8'd87, 8'd126, 8'd87, 8'd106, 8'd82, 8'd110, 8'd134, 8'd129, 8'd161, 8'd75, 8'd130, 8'd50, 8'd64, 8'd127, 8'd142, 8'd155, 8'd117, 8'd175, 8'd152, 8'd160, 8'd148, 8'd132, 8'd109, 8'd130, 8'd86, 8'd71, 8'd91, 8'd134, 8'd134, 8'd93, 8'd159, 8'd166, 8'd105, 8'd140, 8'd105, 8'd138, 8'd73, 8'd133, 8'd55, 8'd55, 8'd78, 8'd110, 8'd66, 8'd120, 8'd127, 8'd101, 8'd115, 8'd106, 8'd76, 8'd136, 8'd99, 8'd128, 8'd34, 8'd143, 8'd141, 8'd116, 8'd87, 8'd165, 8'd129, 8'd100, 8'd103, 8'd146, 8'd96, 8'd154, 8'd78, 8'd105, 8'd39, 8'd63, 8'd45, 8'd90, 8'd123, 8'd135, 8'd98, 8'd167, 8'd150, 8'd93, 8'd120, 8'd71, 8'd123, 8'd96, 8'd32, 8'd116, 8'd121, 8'd94, 8'd104, 8'd91, 8'd101, 8'd123, 8'd127, 8'd118, 8'd153, 8'd63, 8'd111, 8'd59, 8'd134, 8'd131, 8'd82, 8'd85, 8'd58, 8'd112, 8'd79, 8'd129, 8'd94, 8'd141, 8'd173, 8'd109, 8'd100, 8'd128, 8'd103, 8'd124, 8'd68, 8'd148, 8'd156, 8'd166, 8'd126, 8'd136, 8'd180, 8'd163, 8'd145, 8'd134, 8'd77, 8'd137, 8'd58, 8'd79, 8'd107, 8'd92, 8'd86, 8'd139, 8'd60, 8'd144, 8'd182, 8'd140, 8'd87, 8'd80, 8'd146, 8'd56, 8'd127, 8'd75, 8'd116, 8'd156, 8'd133, 8'd102, 8'd138, 8'd116, 8'd156, 8'd152, 8'd142, 8'd134, 8'd70, 8'd131, 8'd56, 8'd146, 8'd69, 8'd95, 8'd101, 8'd80, 8'd133, 8'd189, 8'd170, 8'd97, 8'd92, 8'd154, 8'd136, 8'd63, 8'd70, 8'd56, 8'd85, 8'd121, 8'd108, 8'd141, 8'd139, 8'd153, 8'd173, 8'd172, 8'd104, 8'd131, 8'd104, 8'd147, 8'd111, 8'd94, 8'd127, 8'd161, 8'd122, 8'd129, 8'd141, 8'd130, 8'd141, 8'd136, 8'd102, 8'd79, 8'd132, 8'd161, 8'd158, 8'd34, 8'd44, 8'd86, 8'd103, 8'd56, 8'd75, 8'd145, 8'd176, 8'd153, 8'd183, 8'd158, 8'd174, 8'd157, 8'd112, 8'd108, 8'd71, 8'd173, 8'd146, 8'd102, 8'd132, 8'd113, 8'd141, 8'd139, 8'd145, 8'd95, 8'd138, 8'd143, 8'd187, 8'd137, 8'd139, 8'd110, 8'd140, 8'd64, 8'd102, 8'd89, 8'd103, 8'd106, 8'd136, 8'd176, 8'd119, 8'd147, 8'd95, 8'd166, 8'd109, 8'd110, 8'd85, 8'd144, 8'd136, 8'd142, 8'd181, 8'd122, 8'd129, 8'd116, 8'd132, 8'd157, 8'd206, 8'd203, 8'd170, 8'd151, 8'd169, 8'd110, 8'd168, 8'd77, 8'd140, 8'd156, 8'd137, 8'd95, 8'd105, 8'd171, 8'd150, 8'd174, 8'd129, 8'd168, 8'd186, 8'd128, 8'd120, 8'd182, 8'd100, 8'd153, 8'd157, 8'd133, 8'd118, 8'd169, 8'd142, 8'd155, 8'd148, 8'd182, 8'd165, 8'd162, 8'd144, 8'd155, 8'd102, 8'd76, 8'd120, 8'd90, 8'd174, 8'd163, 8'd186, 8'd181, 8'd161, 8'd101, 8'd116, 8'd179, 8'd159, 8'd135, 8'd124, 8'd150, 8'd118, 8'd165, 8'd115, 8'd160, 8'd195, 8'd130, 8'd171, 8'd168, 8'd155, 8'd183, 8'd161, 8'd97, 8'd159, 8'd137, 8'd170, 8'd127, 8'd103, 8'd178, 8'd150, 8'd95, 8'd110, 8'd149, 8'd171, 8'd170, 8'd96, 8'd111, 8'd110, 8'd136, 8'd165, 8'd142, 8'd92, 8'd102, 8'd109, 8'd152, 8'd167, 8'd135, 8'd107, 8'd89, 8'd156, 8'd126, 8'd190, 8'd141, 8'd117, 8'd133, 8'd144, 8'd141, 8'd108, 8'd168, 8'd118, 8'd122, 8'd95, 8'd135, 8'd129, 8'd118, 8'd142, 8'd174, 8'd179, 8'd138, 8'd146, 8'd141, 8'd125, 8'd149, 8'd109, 8'd156, 8'd113, 8'd97, 8'd114, 8'd153, 8'd108, 8'd118, 8'd145, 8'd83, 8'd147, 8'd180, 8'd137, 8'd157, 8'd131, 8'd166, 8'd161, 8'd149, 8'd139, 8'd114, 8'd152, 8'd180, 8'd138, 8'd83, 8'd99, 8'd116, 8'd97, 8'd144, 8'd124, 8'd125, 8'd157, 8'd142, 8'd145, 8'd96, 8'd98, 8'd131, 8'd86, 8'd88, 8'd117, 8'd164, 8'd114, 8'd102, 8'd110, 8'd159, 8'd144, 8'd100, 8'd110, 8'd90, 8'd168, 8'd146, 8'd156, 8'd103, 8'd90, 8'd76, 8'd120, 8'd90, 8'd115, 8'd110, 8'd105, 8'd108, 8'd83, 8'd98, 8'd64, 8'd124, 8'd82, 8'd59, 8'd125, 8'd76, 8'd117, 8'd121, 8'd72, 8'd67, 8'd102, 8'd147, 8'd113, 8'd94, 8'd145, 8'd156, 8'd102, 8'd119, 8'd138, 8'd111, 8'd109, 8'd146, 8'd111, 8'd113, 8'd125, 8'd139, 8'd165, 8'd128, 8'd153, 8'd76, 8'd85, 8'd64, 8'd75, 8'd153, 8'd75, 8'd127, 8'd103, 8'd82, 8'd91, 8'd98, 8'd144, 8'd95, 8'd112, 8'd106, 8'd125, 8'd168, 8'd85, 8'd118, 8'd61, 8'd61, 8'd109, 8'd131, 8'd67, 8'd73, 8'd83, 8'd63, 8'd145, 8'd40, 8'd42, 8'd94, 8'd84, 8'd14, 8'd29, 8'd74, 8'd104, 8'd79, 8'd97, 8'd106, 8'd132, 8'd153, 8'd133, 8'd75, 8'd169, 8'd83, 8'd168, 8'd135, 8'd85, 8'd115, 8'd145, 8'd65, 8'd150, 8'd135, 8'd53, 8'd95, 8'd72, 8'd56, 8'd43, 8'd57, 8'd110, 8'd59, 8'd117, 8'd48, 8'd130, 8'd75, 8'd87, 8'd92, 8'd102, 8'd80, 8'd136, 8'd115, 8'd71, 8'd111, 8'd73, 8'd77, 8'd104, 8'd138, 8'd157, 8'd126, 8'd160, 8'd114, 8'd118, 8'd96, 8'd99, 8'd130, 8'd151, 8'd141, 8'd100, 8'd151, 8'd145, 8'd82, 8'd159, 8'd99, 8'd137, 8'd81, 8'd90, 8'd104, 8'd80, 8'd160, 8'd113, 8'd74})
) cell_0_89 (
    .clk(clk),
    .input_index(index_0_88_89),
    .input_value(value_0_88_89),
    .input_result(result_0_88_89),
    .input_enable(enable_0_88_89),
    .output_index(index_0_89_90),
    .output_value(value_0_89_90),
    .output_result(result_0_89_90),
    .output_enable(enable_0_89_90)
);

wire [10-1:0] index_0_90_91;
wire [`DATA_WIDTH-1:0] value_0_90_91;
wire [`DATA_WIDTH*4:0] result_0_90_91;
wire enable_0_90_91;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd114, 8'd112, 8'd144, 8'd167, 8'd119, 8'd123, 8'd157, 8'd76, 8'd160, 8'd112, 8'd82, 8'd140, 8'd139, 8'd104, 8'd119, 8'd139, 8'd112, 8'd160, 8'd117, 8'd71, 8'd101, 8'd112, 8'd99, 8'd73, 8'd75, 8'd132, 8'd102, 8'd152, 8'd162, 8'd142, 8'd100, 8'd141, 8'd91, 8'd164, 8'd168, 8'd126, 8'd134, 8'd119, 8'd87, 8'd156, 8'd162, 8'd105, 8'd93, 8'd109, 8'd150, 8'd108, 8'd131, 8'd140, 8'd147, 8'd188, 8'd161, 8'd136, 8'd124, 8'd119, 8'd91, 8'd140, 8'd88, 8'd135, 8'd164, 8'd95, 8'd134, 8'd106, 8'd136, 8'd129, 8'd126, 8'd137, 8'd80, 8'd125, 8'd54, 8'd100, 8'd62, 8'd125, 8'd117, 8'd50, 8'd111, 8'd92, 8'd110, 8'd81, 8'd140, 8'd69, 8'd57, 8'd69, 8'd123, 8'd158, 8'd137, 8'd88, 8'd98, 8'd105, 8'd180, 8'd93, 8'd150, 8'd144, 8'd145, 8'd110, 8'd141, 8'd143, 8'd91, 8'd74, 8'd103, 8'd81, 8'd66, 8'd121, 8'd124, 8'd63, 8'd85, 8'd69, 8'd90, 8'd41, 8'd127, 8'd126, 8'd169, 8'd86, 8'd148, 8'd121, 8'd152, 8'd146, 8'd110, 8'd173, 8'd158, 8'd157, 8'd124, 8'd173, 8'd163, 8'd124, 8'd84, 8'd126, 8'd83, 8'd135, 8'd135, 8'd99, 8'd115, 8'd119, 8'd112, 8'd74, 8'd85, 8'd145, 8'd131, 8'd143, 8'd155, 8'd80, 8'd158, 8'd148, 8'd86, 8'd131, 8'd146, 8'd121, 8'd140, 8'd141, 8'd119, 8'd154, 8'd83, 8'd79, 8'd133, 8'd64, 8'd141, 8'd66, 8'd75, 8'd92, 8'd132, 8'd126, 8'd110, 8'd179, 8'd91, 8'd91, 8'd67, 8'd103, 8'd101, 8'd98, 8'd122, 8'd101, 8'd100, 8'd114, 8'd165, 8'd130, 8'd126, 8'd150, 8'd130, 8'd135, 8'd148, 8'd95, 8'd122, 8'd44, 8'd121, 8'd139, 8'd127, 8'd154, 8'd124, 8'd138, 8'd135, 8'd121, 8'd148, 8'd85, 8'd94, 8'd124, 8'd128, 8'd93, 8'd82, 8'd114, 8'd160, 8'd114, 8'd105, 8'd123, 8'd145, 8'd57, 8'd118, 8'd53, 8'd94, 8'd92, 8'd119, 8'd89, 8'd122, 8'd86, 8'd87, 8'd97, 8'd130, 8'd92, 8'd134, 8'd101, 8'd49, 8'd123, 8'd45, 8'd82, 8'd140, 8'd138, 8'd135, 8'd117, 8'd140, 8'd156, 8'd124, 8'd116, 8'd134, 8'd143, 8'd126, 8'd126, 8'd59, 8'd98, 8'd130, 8'd140, 8'd170, 8'd85, 8'd88, 8'd46, 8'd86, 8'd112, 8'd73, 8'd93, 8'd82, 8'd115, 8'd135, 8'd141, 8'd61, 8'd170, 8'd171, 8'd143, 8'd96, 8'd108, 8'd124, 8'd49, 8'd118, 8'd104, 8'd118, 8'd135, 8'd75, 8'd80, 8'd113, 8'd205, 8'd170, 8'd183, 8'd72, 8'd63, 8'd136, 8'd58, 8'd54, 8'd69, 8'd133, 8'd103, 8'd71, 8'd113, 8'd93, 8'd145, 8'd106, 8'd176, 8'd130, 8'd99, 8'd121, 8'd99, 8'd120, 8'd101, 8'd99, 8'd117, 8'd97, 8'd138, 8'd172, 8'd201, 8'd138, 8'd104, 8'd143, 8'd91, 8'd109, 8'd96, 8'd73, 8'd109, 8'd149, 8'd58, 8'd106, 8'd146, 8'd70, 8'd101, 8'd159, 8'd120, 8'd116, 8'd131, 8'd72, 8'd85, 8'd134, 8'd126, 8'd51, 8'd47, 8'd75, 8'd102, 8'd180, 8'd141, 8'd102, 8'd119, 8'd81, 8'd111, 8'd86, 8'd75, 8'd119, 8'd76, 8'd86, 8'd113, 8'd66, 8'd113, 8'd133, 8'd159, 8'd145, 8'd163, 8'd78, 8'd110, 8'd86, 8'd71, 8'd81, 8'd115, 8'd136, 8'd77, 8'd79, 8'd108, 8'd84, 8'd92, 8'd80, 8'd139, 8'd119, 8'd45, 8'd113, 8'd153, 8'd164, 8'd75, 8'd119, 8'd150, 8'd153, 8'd99, 8'd95, 8'd67, 8'd114, 8'd124, 8'd150, 8'd53, 8'd81, 8'd131, 8'd121, 8'd141, 8'd133, 8'd65, 8'd123, 8'd80, 8'd170, 8'd180, 8'd136, 8'd108, 8'd79, 8'd105, 8'd117, 8'd142, 8'd146, 8'd103, 8'd167, 8'd115, 8'd120, 8'd65, 8'd81, 8'd133, 8'd97, 8'd105, 8'd96, 8'd115, 8'd73, 8'd128, 8'd151, 8'd182, 8'd114, 8'd71, 8'd67, 8'd160, 8'd114, 8'd107, 8'd83, 8'd124, 8'd115, 8'd60, 8'd90, 8'd161, 8'd119, 8'd88, 8'd129, 8'd109, 8'd79, 8'd106, 8'd107, 8'd79, 8'd110, 8'd123, 8'd91, 8'd99, 8'd46, 8'd153, 8'd90, 8'd140, 8'd152, 8'd98, 8'd134, 8'd112, 8'd112, 8'd120, 8'd156, 8'd113, 8'd86, 8'd133, 8'd169, 8'd118, 8'd136, 8'd170, 8'd136, 8'd180, 8'd86, 8'd69, 8'd103, 8'd95, 8'd88, 8'd122, 8'd114, 8'd106, 8'd107, 8'd98, 8'd130, 8'd81, 8'd117, 8'd93, 8'd97, 8'd111, 8'd213, 8'd114, 8'd97, 8'd118, 8'd150, 8'd157, 8'd109, 8'd170, 8'd123, 8'd152, 8'd130, 8'd95, 8'd57, 8'd137, 8'd63, 8'd126, 8'd81, 8'd118, 8'd50, 8'd19, 8'd101, 8'd108, 8'd66, 8'd114, 8'd92, 8'd94, 8'd172, 8'd187, 8'd209, 8'd158, 8'd77, 8'd176, 8'd170, 8'd155, 8'd159, 8'd159, 8'd83, 8'd121, 8'd128, 8'd79, 8'd70, 8'd86, 8'd139, 8'd160, 8'd115, 8'd132, 8'd126, 8'd71, 8'd45, 8'd151, 8'd138, 8'd99, 8'd81, 8'd154, 8'd154, 8'd109, 8'd102, 8'd145, 8'd89, 8'd156, 8'd165, 8'd92, 8'd72, 8'd164, 8'd103, 8'd96, 8'd95, 8'd64, 8'd86, 8'd74, 8'd96, 8'd72, 8'd158, 8'd67, 8'd135, 8'd57, 8'd112, 8'd108, 8'd88, 8'd79, 8'd161, 8'd91, 8'd157, 8'd111, 8'd133, 8'd100, 8'd150, 8'd148, 8'd135, 8'd61, 8'd109, 8'd120, 8'd133, 8'd58, 8'd97, 8'd57, 8'd89, 8'd156, 8'd118, 8'd156, 8'd98, 8'd150, 8'd134, 8'd132, 8'd115, 8'd164, 8'd144, 8'd88, 8'd158, 8'd145, 8'd124, 8'd159, 8'd149, 8'd71, 8'd126, 8'd124, 8'd47, 8'd107, 8'd88, 8'd49, 8'd80, 8'd72, 8'd120, 8'd95, 8'd126, 8'd75, 8'd137, 8'd133, 8'd138, 8'd129, 8'd84, 8'd165, 8'd170, 8'd93, 8'd88, 8'd140, 8'd94, 8'd83, 8'd84, 8'd68, 8'd62, 8'd82, 8'd149, 8'd69, 8'd133, 8'd134, 8'd115, 8'd38, 8'd75, 8'd86, 8'd95, 8'd90, 8'd136, 8'd134, 8'd64, 8'd162, 8'd76, 8'd117, 8'd124, 8'd163, 8'd151, 8'd163, 8'd115, 8'd116, 8'd118, 8'd124, 8'd88, 8'd57, 8'd160, 8'd85, 8'd87, 8'd74, 8'd142, 8'd119, 8'd67, 8'd49, 8'd92, 8'd89, 8'd103, 8'd92, 8'd159, 8'd147, 8'd132, 8'd134, 8'd129, 8'd66, 8'd153, 8'd89, 8'd133, 8'd129, 8'd96, 8'd125, 8'd167, 8'd139, 8'd90, 8'd96, 8'd88, 8'd147, 8'd70, 8'd56, 8'd133, 8'd54, 8'd57, 8'd76, 8'd106, 8'd117, 8'd99, 8'd114, 8'd104, 8'd151, 8'd140, 8'd150, 8'd147, 8'd147, 8'd77, 8'd72, 8'd121, 8'd63, 8'd130, 8'd77, 8'd54, 8'd120, 8'd48, 8'd93, 8'd100, 8'd120, 8'd119, 8'd79, 8'd101, 8'd82, 8'd125, 8'd98, 8'd137, 8'd90, 8'd102, 8'd129, 8'd142, 8'd173, 8'd141, 8'd113, 8'd80, 8'd146, 8'd71, 8'd118, 8'd73, 8'd47, 8'd69, 8'd69, 8'd122, 8'd140, 8'd96, 8'd109, 8'd145, 8'd49, 8'd103, 8'd49, 8'd40, 8'd113, 8'd117, 8'd44, 8'd121, 8'd132, 8'd85, 8'd90, 8'd87, 8'd114, 8'd110, 8'd107, 8'd162, 8'd131, 8'd166, 8'd77, 8'd137, 8'd147, 8'd72, 8'd128, 8'd104, 8'd130, 8'd89, 8'd132, 8'd139, 8'd74, 8'd72, 8'd81, 8'd139, 8'd134, 8'd125, 8'd88, 8'd88, 8'd149, 8'd100, 8'd117, 8'd110, 8'd111, 8'd100, 8'd102, 8'd150, 8'd104, 8'd126, 8'd136, 8'd148, 8'd71, 8'd151, 8'd141, 8'd164, 8'd112, 8'd105, 8'd156, 8'd110, 8'd88, 8'd143, 8'd99, 8'd97, 8'd144, 8'd84, 8'd111, 8'd97, 8'd96, 8'd107, 8'd125, 8'd96, 8'd147, 8'd167, 8'd168})
) cell_0_90 (
    .clk(clk),
    .input_index(index_0_89_90),
    .input_value(value_0_89_90),
    .input_result(result_0_89_90),
    .input_enable(enable_0_89_90),
    .output_index(index_0_90_91),
    .output_value(value_0_90_91),
    .output_result(result_0_90_91),
    .output_enable(enable_0_90_91)
);

wire [10-1:0] index_0_91_92;
wire [`DATA_WIDTH-1:0] value_0_91_92;
wire [`DATA_WIDTH*4:0] result_0_91_92;
wire enable_0_91_92;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd115, 8'd72, 8'd110, 8'd91, 8'd93, 8'd125, 8'd129, 8'd104, 8'd147, 8'd92, 8'd200, 8'd171, 8'd148, 8'd145, 8'd195, 8'd83, 8'd86, 8'd177, 8'd116, 8'd123, 8'd118, 8'd118, 8'd101, 8'd173, 8'd158, 8'd89, 8'd168, 8'd108, 8'd119, 8'd114, 8'd102, 8'd137, 8'd128, 8'd124, 8'd82, 8'd118, 8'd125, 8'd183, 8'd87, 8'd145, 8'd159, 8'd148, 8'd176, 8'd160, 8'd167, 8'd90, 8'd142, 8'd141, 8'd98, 8'd143, 8'd131, 8'd69, 8'd116, 8'd132, 8'd152, 8'd86, 8'd78, 8'd117, 8'd123, 8'd76, 8'd161, 8'd129, 8'd110, 8'd55, 8'd100, 8'd92, 8'd85, 8'd102, 8'd156, 8'd129, 8'd153, 8'd154, 8'd184, 8'd163, 8'd163, 8'd181, 8'd94, 8'd161, 8'd115, 8'd121, 8'd103, 8'd128, 8'd96, 8'd104, 8'd104, 8'd152, 8'd137, 8'd148, 8'd122, 8'd125, 8'd106, 8'd114, 8'd126, 8'd141, 8'd130, 8'd120, 8'd120, 8'd110, 8'd96, 8'd80, 8'd125, 8'd140, 8'd167, 8'd113, 8'd125, 8'd162, 8'd148, 8'd171, 8'd183, 8'd109, 8'd78, 8'd160, 8'd101, 8'd107, 8'd103, 8'd145, 8'd117, 8'd108, 8'd105, 8'd65, 8'd113, 8'd114, 8'd125, 8'd97, 8'd156, 8'd98, 8'd63, 8'd142, 8'd111, 8'd131, 8'd86, 8'd92, 8'd119, 8'd141, 8'd168, 8'd114, 8'd144, 8'd178, 8'd84, 8'd139, 8'd110, 8'd134, 8'd162, 8'd57, 8'd128, 8'd80, 8'd122, 8'd71, 8'd131, 8'd92, 8'd88, 8'd100, 8'd132, 8'd101, 8'd56, 8'd142, 8'd102, 8'd150, 8'd100, 8'd82, 8'd161, 8'd147, 8'd145, 8'd106, 8'd85, 8'd118, 8'd154, 8'd172, 8'd163, 8'd118, 8'd131, 8'd135, 8'd94, 8'd115, 8'd89, 8'd95, 8'd67, 8'd119, 8'd84, 8'd162, 8'd123, 8'd103, 8'd82, 8'd163, 8'd109, 8'd110, 8'd131, 8'd83, 8'd97, 8'd118, 8'd161, 8'd122, 8'd128, 8'd82, 8'd171, 8'd134, 8'd151, 8'd132, 8'd134, 8'd118, 8'd76, 8'd69, 8'd83, 8'd133, 8'd146, 8'd165, 8'd93, 8'd103, 8'd83, 8'd179, 8'd135, 8'd111, 8'd120, 8'd165, 8'd150, 8'd141, 8'd137, 8'd106, 8'd99, 8'd141, 8'd106, 8'd161, 8'd159, 8'd133, 8'd132, 8'd120, 8'd88, 8'd106, 8'd80, 8'd140, 8'd79, 8'd134, 8'd98, 8'd92, 8'd107, 8'd155, 8'd114, 8'd115, 8'd92, 8'd99, 8'd165, 8'd126, 8'd121, 8'd97, 8'd92, 8'd68, 8'd133, 8'd168, 8'd169, 8'd99, 8'd163, 8'd162, 8'd76, 8'd101, 8'd136, 8'd116, 8'd152, 8'd179, 8'd126, 8'd146, 8'd87, 8'd133, 8'd127, 8'd133, 8'd153, 8'd127, 8'd84, 8'd147, 8'd77, 8'd100, 8'd140, 8'd55, 8'd70, 8'd83, 8'd160, 8'd169, 8'd175, 8'd183, 8'd112, 8'd158, 8'd93, 8'd70, 8'd149, 8'd100, 8'd117, 8'd115, 8'd98, 8'd116, 8'd99, 8'd130, 8'd107, 8'd142, 8'd135, 8'd135, 8'd129, 8'd81, 8'd54, 8'd83, 8'd49, 8'd48, 8'd101, 8'd76, 8'd83, 8'd100, 8'd117, 8'd129, 8'd168, 8'd142, 8'd60, 8'd92, 8'd121, 8'd90, 8'd148, 8'd113, 8'd137, 8'd138, 8'd87, 8'd99, 8'd109, 8'd126, 8'd82, 8'd180, 8'd173, 8'd140, 8'd131, 8'd126, 8'd88, 8'd103, 8'd109, 8'd165, 8'd80, 8'd125, 8'd183, 8'd152, 8'd104, 8'd128, 8'd153, 8'd110, 8'd91, 8'd177, 8'd118, 8'd96, 8'd93, 8'd128, 8'd123, 8'd86, 8'd77, 8'd68, 8'd157, 8'd171, 8'd76, 8'd145, 8'd117, 8'd127, 8'd83, 8'd142, 8'd108, 8'd99, 8'd121, 8'd91, 8'd126, 8'd177, 8'd131, 8'd136, 8'd116, 8'd131, 8'd165, 8'd158, 8'd126, 8'd180, 8'd156, 8'd151, 8'd116, 8'd122, 8'd144, 8'd106, 8'd114, 8'd111, 8'd151, 8'd45, 8'd123, 8'd48, 8'd62, 8'd75, 8'd97, 8'd102, 8'd111, 8'd88, 8'd131, 8'd114, 8'd137, 8'd167, 8'd65, 8'd140, 8'd141, 8'd119, 8'd125, 8'd152, 8'd90, 8'd139, 8'd94, 8'd126, 8'd131, 8'd88, 8'd156, 8'd139, 8'd76, 8'd82, 8'd80, 8'd54, 8'd125, 8'd133, 8'd135, 8'd87, 8'd114, 8'd136, 8'd145, 8'd168, 8'd132, 8'd122, 8'd155, 8'd150, 8'd89, 8'd156, 8'd137, 8'd88, 8'd83, 8'd53, 8'd149, 8'd93, 8'd150, 8'd94, 8'd143, 8'd171, 8'd145, 8'd140, 8'd138, 8'd77, 8'd94, 8'd105, 8'd157, 8'd129, 8'd130, 8'd152, 8'd174, 8'd151, 8'd116, 8'd151, 8'd107, 8'd100, 8'd105, 8'd128, 8'd97, 8'd61, 8'd110, 8'd106, 8'd81, 8'd108, 8'd84, 8'd146, 8'd121, 8'd185, 8'd111, 8'd65, 8'd113, 8'd66, 8'd136, 8'd85, 8'd121, 8'd130, 8'd86, 8'd151, 8'd175, 8'd143, 8'd111, 8'd170, 8'd100, 8'd121, 8'd121, 8'd119, 8'd75, 8'd66, 8'd141, 8'd144, 8'd97, 8'd76, 8'd107, 8'd130, 8'd200, 8'd194, 8'd129, 8'd105, 8'd68, 8'd121, 8'd62, 8'd82, 8'd99, 8'd150, 8'd107, 8'd127, 8'd109, 8'd171, 8'd96, 8'd81, 8'd120, 8'd138, 8'd72, 8'd78, 8'd86, 8'd91, 8'd106, 8'd65, 8'd113, 8'd142, 8'd171, 8'd114, 8'd141, 8'd133, 8'd117, 8'd96, 8'd104, 8'd118, 8'd83, 8'd127, 8'd106, 8'd122, 8'd168, 8'd195, 8'd163, 8'd89, 8'd98, 8'd123, 8'd137, 8'd107, 8'd93, 8'd106, 8'd87, 8'd88, 8'd99, 8'd145, 8'd101, 8'd152, 8'd88, 8'd152, 8'd96, 8'd140, 8'd166, 8'd85, 8'd114, 8'd99, 8'd139, 8'd118, 8'd159, 8'd117, 8'd98, 8'd127, 8'd104, 8'd89, 8'd128, 8'd119, 8'd73, 8'd90, 8'd31, 8'd111, 8'd63, 8'd66, 8'd89, 8'd134, 8'd85, 8'd79, 8'd165, 8'd163, 8'd134, 8'd143, 8'd137, 8'd112, 8'd120, 8'd138, 8'd157, 8'd74, 8'd111, 8'd95, 8'd171, 8'd175, 8'd124, 8'd98, 8'd145, 8'd117, 8'd93, 8'd92, 8'd83, 8'd85, 8'd81, 8'd123, 8'd123, 8'd111, 8'd73, 8'd125, 8'd99, 8'd102, 8'd86, 8'd91, 8'd149, 8'd86, 8'd143, 8'd141, 8'd144, 8'd152, 8'd158, 8'd112, 8'd146, 8'd150, 8'd145, 8'd156, 8'd88, 8'd89, 8'd155, 8'd90, 8'd99, 8'd171, 8'd105, 8'd118, 8'd172, 8'd105, 8'd75, 8'd110, 8'd103, 8'd77, 8'd112, 8'd117, 8'd121, 8'd136, 8'd82, 8'd145, 8'd109, 8'd129, 8'd176, 8'd184, 8'd166, 8'd131, 8'd89, 8'd91, 8'd79, 8'd126, 8'd121, 8'd139, 8'd111, 8'd105, 8'd117, 8'd148, 8'd159, 8'd177, 8'd133, 8'd167, 8'd122, 8'd137, 8'd144, 8'd166, 8'd110, 8'd153, 8'd131, 8'd99, 8'd92, 8'd142, 8'd96, 8'd153, 8'd186, 8'd147, 8'd99, 8'd142, 8'd152, 8'd150, 8'd104, 8'd135, 8'd95, 8'd152, 8'd142, 8'd158, 8'd143, 8'd173, 8'd118, 8'd141, 8'd134, 8'd122, 8'd166, 8'd154, 8'd137, 8'd195, 8'd131, 8'd152, 8'd150, 8'd142, 8'd176, 8'd143, 8'd169, 8'd111, 8'd92, 8'd105, 8'd95, 8'd169, 8'd82, 8'd89, 8'd135, 8'd158, 8'd134, 8'd104, 8'd101, 8'd98, 8'd173, 8'd192, 8'd157, 8'd126, 8'd137, 8'd198, 8'd180, 8'd137, 8'd118, 8'd152, 8'd177, 8'd158, 8'd134, 8'd125, 8'd150, 8'd80, 8'd163, 8'd169, 8'd145, 8'd103, 8'd90, 8'd75, 8'd103, 8'd82, 8'd134, 8'd181, 8'd87, 8'd121, 8'd97, 8'd151, 8'd92, 8'd154, 8'd166, 8'd120, 8'd140, 8'd183, 8'd111, 8'd125, 8'd107, 8'd102, 8'd152, 8'd164, 8'd167, 8'd137, 8'd159, 8'd104, 8'd71, 8'd140, 8'd155, 8'd105, 8'd102, 8'd75, 8'd149, 8'd161, 8'd84, 8'd97, 8'd169, 8'd146, 8'd80, 8'd148, 8'd126, 8'd71, 8'd83, 8'd78, 8'd81, 8'd140, 8'd80, 8'd142, 8'd164, 8'd144, 8'd125, 8'd110, 8'd118, 8'd124, 8'd138, 8'd134})
) cell_0_91 (
    .clk(clk),
    .input_index(index_0_90_91),
    .input_value(value_0_90_91),
    .input_result(result_0_90_91),
    .input_enable(enable_0_90_91),
    .output_index(index_0_91_92),
    .output_value(value_0_91_92),
    .output_result(result_0_91_92),
    .output_enable(enable_0_91_92)
);

wire [10-1:0] index_0_92_93;
wire [`DATA_WIDTH-1:0] value_0_92_93;
wire [`DATA_WIDTH*4:0] result_0_92_93;
wire enable_0_92_93;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd132, 8'd76, 8'd97, 8'd169, 8'd59, 8'd128, 8'd147, 8'd119, 8'd126, 8'd119, 8'd76, 8'd80, 8'd57, 8'd66, 8'd92, 8'd88, 8'd112, 8'd84, 8'd102, 8'd139, 8'd144, 8'd85, 8'd148, 8'd93, 8'd135, 8'd117, 8'd109, 8'd97, 8'd118, 8'd74, 8'd95, 8'd116, 8'd139, 8'd67, 8'd104, 8'd127, 8'd70, 8'd67, 8'd149, 8'd76, 8'd144, 8'd119, 8'd124, 8'd79, 8'd151, 8'd67, 8'd75, 8'd126, 8'd140, 8'd138, 8'd135, 8'd166, 8'd167, 8'd81, 8'd157, 8'd123, 8'd152, 8'd91, 8'd87, 8'd96, 8'd119, 8'd135, 8'd110, 8'd188, 8'd166, 8'd108, 8'd86, 8'd125, 8'd94, 8'd113, 8'd106, 8'd126, 8'd76, 8'd72, 8'd89, 8'd105, 8'd84, 8'd86, 8'd93, 8'd148, 8'd148, 8'd162, 8'd90, 8'd139, 8'd117, 8'd115, 8'd128, 8'd161, 8'd209, 8'd153, 8'd198, 8'd152, 8'd121, 8'd151, 8'd147, 8'd151, 8'd142, 8'd143, 8'd77, 8'd60, 8'd57, 8'd149, 8'd155, 8'd152, 8'd65, 8'd87, 8'd106, 8'd113, 8'd74, 8'd129, 8'd120, 8'd148, 8'd76, 8'd168, 8'd160, 8'd163, 8'd170, 8'd161, 8'd137, 8'd172, 8'd120, 8'd144, 8'd138, 8'd133, 8'd162, 8'd72, 8'd84, 8'd75, 8'd87, 8'd121, 8'd94, 8'd154, 8'd77, 8'd79, 8'd100, 8'd144, 8'd101, 8'd158, 8'd169, 8'd147, 8'd109, 8'd104, 8'd152, 8'd163, 8'd132, 8'd154, 8'd120, 8'd175, 8'd103, 8'd169, 8'd86, 8'd83, 8'd140, 8'd144, 8'd114, 8'd86, 8'd168, 8'd158, 8'd139, 8'd157, 8'd100, 8'd199, 8'd131, 8'd116, 8'd145, 8'd114, 8'd110, 8'd163, 8'd131, 8'd101, 8'd179, 8'd122, 8'd104, 8'd101, 8'd189, 8'd195, 8'd176, 8'd92, 8'd97, 8'd93, 8'd83, 8'd63, 8'd65, 8'd78, 8'd80, 8'd112, 8'd122, 8'd170, 8'd175, 8'd125, 8'd130, 8'd170, 8'd212, 8'd131, 8'd82, 8'd83, 8'd161, 8'd115, 8'd192, 8'd132, 8'd186, 8'd193, 8'd115, 8'd155, 8'd157, 8'd153, 8'd175, 8'd154, 8'd71, 8'd129, 8'd146, 8'd134, 8'd143, 8'd126, 8'd125, 8'd126, 8'd165, 8'd201, 8'd154, 8'd190, 8'd150, 8'd159, 8'd159, 8'd137, 8'd117, 8'd139, 8'd182, 8'd145, 8'd175, 8'd113, 8'd129, 8'd120, 8'd106, 8'd165, 8'd124, 8'd84, 8'd148, 8'd81, 8'd137, 8'd124, 8'd95, 8'd70, 8'd145, 8'd147, 8'd173, 8'd140, 8'd160, 8'd184, 8'd171, 8'd160, 8'd113, 8'd115, 8'd135, 8'd111, 8'd101, 8'd102, 8'd157, 8'd153, 8'd102, 8'd147, 8'd157, 8'd115, 8'd155, 8'd83, 8'd131, 8'd85, 8'd140, 8'd101, 8'd61, 8'd52, 8'd119, 8'd119, 8'd135, 8'd165, 8'd137, 8'd158, 8'd126, 8'd113, 8'd163, 8'd155, 8'd163, 8'd164, 8'd167, 8'd102, 8'd125, 8'd117, 8'd156, 8'd77, 8'd70, 8'd101, 8'd66, 8'd163, 8'd89, 8'd127, 8'd137, 8'd79, 8'd51, 8'd74, 8'd118, 8'd80, 8'd153, 8'd110, 8'd169, 8'd153, 8'd183, 8'd147, 8'd139, 8'd146, 8'd148, 8'd136, 8'd138, 8'd145, 8'd87, 8'd146, 8'd88, 8'd148, 8'd60, 8'd97, 8'd73, 8'd111, 8'd133, 8'd150, 8'd181, 8'd137, 8'd134, 8'd105, 8'd129, 8'd127, 8'd91, 8'd94, 8'd166, 8'd122, 8'd161, 8'd81, 8'd126, 8'd157, 8'd95, 8'd203, 8'd157, 8'd80, 8'd44, 8'd53, 8'd72, 8'd97, 8'd109, 8'd134, 8'd79, 8'd79, 8'd142, 8'd169, 8'd170, 8'd153, 8'd145, 8'd116, 8'd168, 8'd111, 8'd81, 8'd110, 8'd112, 8'd98, 8'd130, 8'd94, 8'd121, 8'd169, 8'd139, 8'd124, 8'd97, 8'd72, 8'd53, 8'd58, 8'd64, 8'd114, 8'd119, 8'd79, 8'd117, 8'd164, 8'd161, 8'd150, 8'd170, 8'd144, 8'd163, 8'd144, 8'd101, 8'd115, 8'd95, 8'd97, 8'd81, 8'd119, 8'd75, 8'd83, 8'd77, 8'd98, 8'd149, 8'd166, 8'd168, 8'd30, 8'd35, 8'd38, 8'd100, 8'd113, 8'd120, 8'd105, 8'd80, 8'd96, 8'd134, 8'd165, 8'd176, 8'd184, 8'd114, 8'd61, 8'd130, 8'd108, 8'd54, 8'd113, 8'd121, 8'd138, 8'd109, 8'd107, 8'd122, 8'd111, 8'd146, 8'd146, 8'd119, 8'd112, 8'd78, 8'd31, 8'd147, 8'd92, 8'd110, 8'd109, 8'd108, 8'd121, 8'd176, 8'd141, 8'd153, 8'd78, 8'd114, 8'd64, 8'd110, 8'd112, 8'd124, 8'd122, 8'd109, 8'd114, 8'd93, 8'd78, 8'd107, 8'd164, 8'd121, 8'd167, 8'd139, 8'd113, 8'd119, 8'd130, 8'd45, 8'd108, 8'd69, 8'd121, 8'd110, 8'd113, 8'd181, 8'd101, 8'd117, 8'd115, 8'd105, 8'd146, 8'd115, 8'd122, 8'd128, 8'd78, 8'd146, 8'd84, 8'd110, 8'd63, 8'd75, 8'd131, 8'd167, 8'd109, 8'd198, 8'd163, 8'd75, 8'd110, 8'd140, 8'd72, 8'd106, 8'd136, 8'd76, 8'd119, 8'd112, 8'd135, 8'd105, 8'd67, 8'd144, 8'd91, 8'd61, 8'd109, 8'd61, 8'd144, 8'd149, 8'd91, 8'd131, 8'd127, 8'd88, 8'd97, 8'd136, 8'd143, 8'd163, 8'd100, 8'd92, 8'd73, 8'd95, 8'd104, 8'd152, 8'd88, 8'd88, 8'd86, 8'd141, 8'd122, 8'd137, 8'd157, 8'd125, 8'd109, 8'd66, 8'd124, 8'd84, 8'd130, 8'd104, 8'd97, 8'd55, 8'd120, 8'd135, 8'd158, 8'd128, 8'd167, 8'd185, 8'd87, 8'd96, 8'd134, 8'd123, 8'd96, 8'd92, 8'd125, 8'd83, 8'd91, 8'd119, 8'd111, 8'd159, 8'd82, 8'd55, 8'd124, 8'd128, 8'd137, 8'd117, 8'd71, 8'd64, 8'd127, 8'd99, 8'd93, 8'd122, 8'd141, 8'd82, 8'd129, 8'd119, 8'd154, 8'd100, 8'd143, 8'd119, 8'd88, 8'd155, 8'd104, 8'd165, 8'd99, 8'd120, 8'd184, 8'd133, 8'd91, 8'd125, 8'd62, 8'd114, 8'd108, 8'd43, 8'd63, 8'd81, 8'd124, 8'd95, 8'd78, 8'd100, 8'd110, 8'd110, 8'd123, 8'd92, 8'd144, 8'd65, 8'd79, 8'd144, 8'd99, 8'd103, 8'd112, 8'd111, 8'd95, 8'd173, 8'd152, 8'd146, 8'd97, 8'd110, 8'd62, 8'd106, 8'd107, 8'd72, 8'd131, 8'd142, 8'd147, 8'd106, 8'd60, 8'd171, 8'd127, 8'd84, 8'd150, 8'd72, 8'd94, 8'd129, 8'd49, 8'd93, 8'd162, 8'd80, 8'd78, 8'd138, 8'd96, 8'd104, 8'd126, 8'd118, 8'd120, 8'd189, 8'd96, 8'd67, 8'd82, 8'd69, 8'd99, 8'd157, 8'd166, 8'd173, 8'd113, 8'd112, 8'd133, 8'd114, 8'd142, 8'd100, 8'd117, 8'd127, 8'd103, 8'd122, 8'd106, 8'd56, 8'd96, 8'd112, 8'd163, 8'd117, 8'd164, 8'd130, 8'd163, 8'd190, 8'd170, 8'd179, 8'd75, 8'd138, 8'd149, 8'd114, 8'd125, 8'd149, 8'd134, 8'd82, 8'd72, 8'd73, 8'd92, 8'd88, 8'd125, 8'd95, 8'd99, 8'd81, 8'd68, 8'd101, 8'd90, 8'd104, 8'd90, 8'd108, 8'd141, 8'd78, 8'd111, 8'd111, 8'd116, 8'd108, 8'd72, 8'd135, 8'd141, 8'd117, 8'd162, 8'd103, 8'd140, 8'd77, 8'd82, 8'd128, 8'd74, 8'd124, 8'd154, 8'd95, 8'd58, 8'd133, 8'd84, 8'd59, 8'd65, 8'd127, 8'd106, 8'd98, 8'd144, 8'd64, 8'd101, 8'd97, 8'd105, 8'd60, 8'd47, 8'd115, 8'd53, 8'd117, 8'd98, 8'd125, 8'd167, 8'd91, 8'd79, 8'd143, 8'd134, 8'd157, 8'd146, 8'd107, 8'd106, 8'd63, 8'd135, 8'd79, 8'd99, 8'd115, 8'd76, 8'd138, 8'd126, 8'd74, 8'd119, 8'd60, 8'd125, 8'd61, 8'd64, 8'd83, 8'd84, 8'd154, 8'd81, 8'd94, 8'd167, 8'd138, 8'd127, 8'd87, 8'd144, 8'd83, 8'd105, 8'd155, 8'd125, 8'd159, 8'd74, 8'd103, 8'd124, 8'd143, 8'd160, 8'd163, 8'd152, 8'd86, 8'd128, 8'd128, 8'd74, 8'd167, 8'd145, 8'd81, 8'd115, 8'd98, 8'd127, 8'd108, 8'd70, 8'd86, 8'd72})
) cell_0_92 (
    .clk(clk),
    .input_index(index_0_91_92),
    .input_value(value_0_91_92),
    .input_result(result_0_91_92),
    .input_enable(enable_0_91_92),
    .output_index(index_0_92_93),
    .output_value(value_0_92_93),
    .output_result(result_0_92_93),
    .output_enable(enable_0_92_93)
);

wire [10-1:0] index_0_93_94;
wire [`DATA_WIDTH-1:0] value_0_93_94;
wire [`DATA_WIDTH*4:0] result_0_93_94;
wire enable_0_93_94;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd83, 8'd126, 8'd72, 8'd123, 8'd84, 8'd80, 8'd137, 8'd155, 8'd101, 8'd79, 8'd112, 8'd103, 8'd82, 8'd124, 8'd119, 8'd163, 8'd122, 8'd96, 8'd136, 8'd88, 8'd134, 8'd107, 8'd84, 8'd97, 8'd78, 8'd109, 8'd164, 8'd93, 8'd85, 8'd146, 8'd78, 8'd141, 8'd91, 8'd119, 8'd161, 8'd159, 8'd101, 8'd130, 8'd92, 8'd104, 8'd183, 8'd160, 8'd167, 8'd114, 8'd149, 8'd136, 8'd169, 8'd107, 8'd109, 8'd107, 8'd81, 8'd171, 8'd153, 8'd141, 8'd118, 8'd72, 8'd170, 8'd71, 8'd85, 8'd79, 8'd90, 8'd92, 8'd128, 8'd178, 8'd139, 8'd170, 8'd158, 8'd139, 8'd139, 8'd115, 8'd192, 8'd219, 8'd175, 8'd188, 8'd115, 8'd161, 8'd95, 8'd181, 8'd113, 8'd83, 8'd135, 8'd110, 8'd162, 8'd75, 8'd75, 8'd83, 8'd142, 8'd77, 8'd168, 8'd154, 8'd131, 8'd150, 8'd125, 8'd147, 8'd176, 8'd193, 8'd155, 8'd113, 8'd127, 8'd172, 8'd167, 8'd200, 8'd154, 8'd195, 8'd173, 8'd101, 8'd135, 8'd151, 8'd86, 8'd165, 8'd133, 8'd77, 8'd82, 8'd100, 8'd139, 8'd95, 8'd83, 8'd84, 8'd86, 8'd128, 8'd140, 8'd136, 8'd177, 8'd174, 8'd142, 8'd171, 8'd179, 8'd125, 8'd151, 8'd163, 8'd131, 8'd164, 8'd105, 8'd171, 8'd97, 8'd69, 8'd156, 8'd94, 8'd88, 8'd156, 8'd82, 8'd151, 8'd157, 8'd85, 8'd130, 8'd130, 8'd155, 8'd97, 8'd160, 8'd85, 8'd167, 8'd167, 8'd144, 8'd133, 8'd174, 8'd104, 8'd164, 8'd94, 8'd133, 8'd141, 8'd151, 8'd122, 8'd96, 8'd70, 8'd169, 8'd105, 8'd143, 8'd123, 8'd69, 8'd87, 8'd84, 8'd96, 8'd123, 8'd123, 8'd91, 8'd105, 8'd100, 8'd168, 8'd99, 8'd154, 8'd163, 8'd90, 8'd63, 8'd143, 8'd68, 8'd104, 8'd137, 8'd167, 8'd170, 8'd192, 8'd167, 8'd140, 8'd123, 8'd130, 8'd114, 8'd112, 8'd167, 8'd72, 8'd81, 8'd129, 8'd141, 8'd144, 8'd90, 8'd168, 8'd143, 8'd99, 8'd81, 8'd63, 8'd149, 8'd129, 8'd75, 8'd95, 8'd101, 8'd142, 8'd77, 8'd90, 8'd154, 8'd117, 8'd146, 8'd179, 8'd98, 8'd102, 8'd140, 8'd96, 8'd123, 8'd64, 8'd79, 8'd102, 8'd164, 8'd102, 8'd94, 8'd121, 8'd124, 8'd96, 8'd134, 8'd76, 8'd145, 8'd112, 8'd100, 8'd54, 8'd88, 8'd68, 8'd87, 8'd133, 8'd114, 8'd147, 8'd194, 8'd177, 8'd123, 8'd137, 8'd98, 8'd95, 8'd150, 8'd147, 8'd65, 8'd62, 8'd90, 8'd140, 8'd154, 8'd122, 8'd109, 8'd158, 8'd156, 8'd100, 8'd120, 8'd60, 8'd38, 8'd64, 8'd63, 8'd101, 8'd154, 8'd98, 8'd140, 8'd109, 8'd149, 8'd121, 8'd198, 8'd138, 8'd107, 8'd117, 8'd81, 8'd161, 8'd84, 8'd126, 8'd80, 8'd128, 8'd96, 8'd141, 8'd148, 8'd107, 8'd122, 8'd120, 8'd151, 8'd144, 8'd108, 8'd104, 8'd72, 8'd48, 8'd67, 8'd104, 8'd81, 8'd61, 8'd143, 8'd117, 8'd183, 8'd148, 8'd165, 8'd166, 8'd87, 8'd171, 8'd111, 8'd154, 8'd144, 8'd156, 8'd119, 8'd100, 8'd99, 8'd160, 8'd113, 8'd145, 8'd76, 8'd160, 8'd131, 8'd119, 8'd132, 8'd86, 8'd87, 8'd137, 8'd95, 8'd100, 8'd82, 8'd134, 8'd144, 8'd109, 8'd121, 8'd103, 8'd142, 8'd165, 8'd104, 8'd89, 8'd73, 8'd70, 8'd61, 8'd152, 8'd124, 8'd173, 8'd107, 8'd128, 8'd98, 8'd98, 8'd148, 8'd97, 8'd113, 8'd111, 8'd124, 8'd62, 8'd117, 8'd76, 8'd144, 8'd86, 8'd157, 8'd150, 8'd175, 8'd139, 8'd93, 8'd119, 8'd97, 8'd135, 8'd73, 8'd66, 8'd99, 8'd133, 8'd110, 8'd106, 8'd163, 8'd186, 8'd119, 8'd173, 8'd112, 8'd162, 8'd63, 8'd106, 8'd133, 8'd99, 8'd90, 8'd92, 8'd63, 8'd159, 8'd100, 8'd70, 8'd159, 8'd92, 8'd87, 8'd101, 8'd139, 8'd127, 8'd55, 8'd99, 8'd86, 8'd143, 8'd188, 8'd120, 8'd168, 8'd184, 8'd180, 8'd116, 8'd99, 8'd165, 8'd61, 8'd64, 8'd98, 8'd152, 8'd115, 8'd143, 8'd133, 8'd153, 8'd88, 8'd140, 8'd81, 8'd137, 8'd137, 8'd139, 8'd106, 8'd118, 8'd183, 8'd117, 8'd100, 8'd141, 8'd130, 8'd195, 8'd195, 8'd158, 8'd150, 8'd128, 8'd102, 8'd87, 8'd137, 8'd99, 8'd85, 8'd116, 8'd130, 8'd69, 8'd124, 8'd173, 8'd82, 8'd75, 8'd77, 8'd75, 8'd129, 8'd156, 8'd142, 8'd166, 8'd134, 8'd135, 8'd137, 8'd137, 8'd168, 8'd137, 8'd152, 8'd179, 8'd185, 8'd144, 8'd154, 8'd90, 8'd160, 8'd150, 8'd115, 8'd109, 8'd138, 8'd98, 8'd186, 8'd117, 8'd83, 8'd77, 8'd140, 8'd110, 8'd148, 8'd90, 8'd56, 8'd149, 8'd149, 8'd173, 8'd160, 8'd164, 8'd189, 8'd170, 8'd183, 8'd125, 8'd157, 8'd145, 8'd122, 8'd132, 8'd160, 8'd141, 8'd87, 8'd89, 8'd146, 8'd121, 8'd180, 8'd173, 8'd169, 8'd120, 8'd143, 8'd111, 8'd84, 8'd140, 8'd153, 8'd79, 8'd149, 8'd152, 8'd190, 8'd177, 8'd155, 8'd139, 8'd119, 8'd132, 8'd122, 8'd160, 8'd106, 8'd114, 8'd139, 8'd171, 8'd173, 8'd130, 8'd166, 8'd128, 8'd116, 8'd158, 8'd144, 8'd61, 8'd76, 8'd123, 8'd165, 8'd130, 8'd86, 8'd103, 8'd154, 8'd102, 8'd114, 8'd127, 8'd200, 8'd125, 8'd190, 8'd183, 8'd137, 8'd160, 8'd135, 8'd121, 8'd156, 8'd159, 8'd108, 8'd199, 8'd186, 8'd115, 8'd152, 8'd184, 8'd122, 8'd92, 8'd122, 8'd157, 8'd89, 8'd156, 8'd77, 8'd83, 8'd60, 8'd78, 8'd164, 8'd158, 8'd186, 8'd122, 8'd112, 8'd152, 8'd171, 8'd203, 8'd140, 8'd152, 8'd144, 8'd132, 8'd148, 8'd147, 8'd115, 8'd98, 8'd110, 8'd115, 8'd140, 8'd135, 8'd118, 8'd121, 8'd113, 8'd70, 8'd128, 8'd61, 8'd75, 8'd28, 8'd142, 8'd153, 8'd101, 8'd128, 8'd123, 8'd194, 8'd134, 8'd182, 8'd126, 8'd163, 8'd148, 8'd151, 8'd198, 8'd148, 8'd128, 8'd101, 8'd172, 8'd167, 8'd126, 8'd152, 8'd119, 8'd160, 8'd84, 8'd88, 8'd96, 8'd83, 8'd58, 8'd34, 8'd76, 8'd58, 8'd76, 8'd119, 8'd65, 8'd136, 8'd86, 8'd124, 8'd192, 8'd129, 8'd151, 8'd130, 8'd100, 8'd143, 8'd90, 8'd112, 8'd170, 8'd178, 8'd167, 8'd157, 8'd122, 8'd162, 8'd72, 8'd110, 8'd69, 8'd30, 8'd91, 8'd88, 8'd92, 8'd94, 8'd60, 8'd110, 8'd37, 8'd119, 8'd130, 8'd102, 8'd85, 8'd113, 8'd100, 8'd179, 8'd119, 8'd91, 8'd102, 8'd84, 8'd135, 8'd146, 8'd165, 8'd127, 8'd93, 8'd118, 8'd145, 8'd151, 8'd93, 8'd123, 8'd103, 8'd45, 8'd54, 8'd44, 8'd51, 8'd106, 8'd57, 8'd132, 8'd91, 8'd74, 8'd141, 8'd70, 8'd155, 8'd100, 8'd102, 8'd135, 8'd105, 8'd104, 8'd122, 8'd96, 8'd117, 8'd103, 8'd125, 8'd166, 8'd161, 8'd130, 8'd167, 8'd79, 8'd51, 8'd104, 8'd109, 8'd61, 8'd49, 8'd90, 8'd126, 8'd63, 8'd114, 8'd111, 8'd76, 8'd98, 8'd63, 8'd111, 8'd93, 8'd65, 8'd128, 8'd89, 8'd157, 8'd107, 8'd111, 8'd141, 8'd111, 8'd141, 8'd159, 8'd102, 8'd166, 8'd126, 8'd148, 8'd165, 8'd154, 8'd136, 8'd113, 8'd137, 8'd164, 8'd124, 8'd100, 8'd164, 8'd126, 8'd80, 8'd90, 8'd146, 8'd132, 8'd140, 8'd144, 8'd107, 8'd99, 8'd122, 8'd96, 8'd127, 8'd76, 8'd150, 8'd158, 8'd137, 8'd80, 8'd74, 8'd138, 8'd123, 8'd162, 8'd168, 8'd83, 8'd161, 8'd85, 8'd160, 8'd161, 8'd149, 8'd157, 8'd117, 8'd119, 8'd147, 8'd114, 8'd123, 8'd170, 8'd70, 8'd132, 8'd125, 8'd126, 8'd90, 8'd70, 8'd159})
) cell_0_93 (
    .clk(clk),
    .input_index(index_0_92_93),
    .input_value(value_0_92_93),
    .input_result(result_0_92_93),
    .input_enable(enable_0_92_93),
    .output_index(index_0_93_94),
    .output_value(value_0_93_94),
    .output_result(result_0_93_94),
    .output_enable(enable_0_93_94)
);

wire [10-1:0] index_0_94_95;
wire [`DATA_WIDTH-1:0] value_0_94_95;
wire [`DATA_WIDTH*4:0] result_0_94_95;
wire enable_0_94_95;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd128, 8'd119, 8'd153, 8'd101, 8'd133, 8'd135, 8'd121, 8'd92, 8'd113, 8'd107, 8'd92, 8'd106, 8'd117, 8'd107, 8'd100, 8'd71, 8'd127, 8'd143, 8'd155, 8'd120, 8'd170, 8'd88, 8'd74, 8'd162, 8'd88, 8'd159, 8'd128, 8'd112, 8'd89, 8'd158, 8'd93, 8'd143, 8'd87, 8'd156, 8'd150, 8'd77, 8'd91, 8'd137, 8'd92, 8'd156, 8'd121, 8'd144, 8'd144, 8'd150, 8'd145, 8'd80, 8'd101, 8'd116, 8'd108, 8'd97, 8'd129, 8'd124, 8'd122, 8'd130, 8'd121, 8'd153, 8'd85, 8'd115, 8'd111, 8'd100, 8'd161, 8'd104, 8'd136, 8'd122, 8'd163, 8'd97, 8'd79, 8'd108, 8'd124, 8'd74, 8'd155, 8'd124, 8'd142, 8'd109, 8'd100, 8'd118, 8'd128, 8'd97, 8'd142, 8'd89, 8'd134, 8'd173, 8'd74, 8'd101, 8'd105, 8'd102, 8'd157, 8'd82, 8'd81, 8'd142, 8'd101, 8'd148, 8'd91, 8'd112, 8'd137, 8'd165, 8'd140, 8'd138, 8'd118, 8'd192, 8'd114, 8'd180, 8'd136, 8'd110, 8'd162, 8'd91, 8'd119, 8'd83, 8'd126, 8'd144, 8'd116, 8'd159, 8'd94, 8'd164, 8'd99, 8'd105, 8'd128, 8'd103, 8'd117, 8'd122, 8'd122, 8'd143, 8'd120, 8'd116, 8'd118, 8'd154, 8'd143, 8'd189, 8'd145, 8'd96, 8'd115, 8'd92, 8'd128, 8'd154, 8'd81, 8'd171, 8'd152, 8'd175, 8'd129, 8'd129, 8'd163, 8'd144, 8'd156, 8'd108, 8'd129, 8'd155, 8'd168, 8'd132, 8'd85, 8'd172, 8'd168, 8'd151, 8'd82, 8'd181, 8'd107, 8'd154, 8'd170, 8'd82, 8'd77, 8'd153, 8'd106, 8'd120, 8'd163, 8'd93, 8'd93, 8'd90, 8'd155, 8'd96, 8'd150, 8'd96, 8'd157, 8'd138, 8'd69, 8'd124, 8'd138, 8'd104, 8'd116, 8'd100, 8'd130, 8'd169, 8'd159, 8'd101, 8'd103, 8'd150, 8'd84, 8'd137, 8'd166, 8'd91, 8'd185, 8'd132, 8'd168, 8'd104, 8'd180, 8'd166, 8'd85, 8'd112, 8'd88, 8'd138, 8'd85, 8'd148, 8'd99, 8'd162, 8'd182, 8'd148, 8'd94, 8'd117, 8'd157, 8'd158, 8'd118, 8'd145, 8'd92, 8'd130, 8'd113, 8'd147, 8'd122, 8'd185, 8'd134, 8'd170, 8'd159, 8'd139, 8'd194, 8'd170, 8'd135, 8'd132, 8'd78, 8'd134, 8'd95, 8'd104, 8'd149, 8'd142, 8'd127, 8'd175, 8'd176, 8'd118, 8'd162, 8'd166, 8'd76, 8'd76, 8'd146, 8'd88, 8'd110, 8'd99, 8'd141, 8'd133, 8'd140, 8'd142, 8'd112, 8'd173, 8'd153, 8'd140, 8'd167, 8'd133, 8'd60, 8'd136, 8'd119, 8'd132, 8'd180, 8'd113, 8'd184, 8'd169, 8'd158, 8'd144, 8'd146, 8'd89, 8'd63, 8'd95, 8'd133, 8'd55, 8'd109, 8'd87, 8'd115, 8'd108, 8'd131, 8'd127, 8'd123, 8'd128, 8'd156, 8'd126, 8'd104, 8'd86, 8'd146, 8'd84, 8'd93, 8'd90, 8'd152, 8'd126, 8'd118, 8'd76, 8'd172, 8'd112, 8'd127, 8'd135, 8'd48, 8'd34, 8'd68, 8'd92, 8'd94, 8'd105, 8'd154, 8'd89, 8'd107, 8'd89, 8'd153, 8'd164, 8'd131, 8'd126, 8'd125, 8'd148, 8'd106, 8'd120, 8'd100, 8'd101, 8'd187, 8'd147, 8'd106, 8'd102, 8'd99, 8'd133, 8'd148, 8'd111, 8'd61, 8'd105, 8'd119, 8'd150, 8'd162, 8'd143, 8'd151, 8'd101, 8'd99, 8'd78, 8'd98, 8'd169, 8'd92, 8'd155, 8'd134, 8'd164, 8'd86, 8'd88, 8'd132, 8'd200, 8'd97, 8'd78, 8'd120, 8'd156, 8'd99, 8'd105, 8'd100, 8'd71, 8'd104, 8'd96, 8'd188, 8'd104, 8'd97, 8'd137, 8'd117, 8'd161, 8'd94, 8'd64, 8'd98, 8'd143, 8'd102, 8'd166, 8'd80, 8'd115, 8'd141, 8'd100, 8'd135, 8'd154, 8'd117, 8'd83, 8'd124, 8'd84, 8'd105, 8'd112, 8'd71, 8'd123, 8'd93, 8'd181, 8'd106, 8'd108, 8'd119, 8'd64, 8'd73, 8'd87, 8'd84, 8'd136, 8'd74, 8'd78, 8'd145, 8'd94, 8'd153, 8'd76, 8'd142, 8'd166, 8'd111, 8'd143, 8'd94, 8'd159, 8'd85, 8'd104, 8'd75, 8'd125, 8'd113, 8'd92, 8'd90, 8'd121, 8'd142, 8'd131, 8'd105, 8'd148, 8'd84, 8'd125, 8'd126, 8'd127, 8'd49, 8'd91, 8'd124, 8'd115, 8'd75, 8'd90, 8'd148, 8'd95, 8'd183, 8'd126, 8'd169, 8'd97, 8'd161, 8'd124, 8'd108, 8'd139, 8'd88, 8'd81, 8'd147, 8'd124, 8'd135, 8'd155, 8'd139, 8'd75, 8'd69, 8'd67, 8'd71, 8'd86, 8'd70, 8'd71, 8'd95, 8'd159, 8'd139, 8'd123, 8'd82, 8'd161, 8'd167, 8'd198, 8'd170, 8'd172, 8'd108, 8'd156, 8'd95, 8'd143, 8'd81, 8'd138, 8'd106, 8'd117, 8'd154, 8'd114, 8'd94, 8'd62, 8'd109, 8'd89, 8'd70, 8'd94, 8'd151, 8'd83, 8'd171, 8'd162, 8'd161, 8'd159, 8'd175, 8'd165, 8'd97, 8'd186, 8'd156, 8'd150, 8'd160, 8'd167, 8'd129, 8'd151, 8'd116, 8'd91, 8'd160, 8'd116, 8'd86, 8'd61, 8'd83, 8'd87, 8'd72, 8'd108, 8'd131, 8'd104, 8'd118, 8'd118, 8'd130, 8'd113, 8'd159, 8'd91, 8'd75, 8'd175, 8'd129, 8'd113, 8'd164, 8'd100, 8'd163, 8'd128, 8'd112, 8'd107, 8'd130, 8'd128, 8'd159, 8'd108, 8'd83, 8'd154, 8'd113, 8'd152, 8'd118, 8'd127, 8'd152, 8'd139, 8'd96, 8'd152, 8'd158, 8'd155, 8'd96, 8'd152, 8'd88, 8'd138, 8'd97, 8'd82, 8'd95, 8'd88, 8'd133, 8'd163, 8'd138, 8'd162, 8'd133, 8'd101, 8'd159, 8'd192, 8'd113, 8'd133, 8'd136, 8'd157, 8'd140, 8'd78, 8'd161, 8'd135, 8'd107, 8'd115, 8'd147, 8'd69, 8'd115, 8'd111, 8'd136, 8'd156, 8'd74, 8'd96, 8'd159, 8'd124, 8'd105, 8'd153, 8'd165, 8'd152, 8'd170, 8'd182, 8'd137, 8'd156, 8'd120, 8'd102, 8'd119, 8'd150, 8'd135, 8'd90, 8'd147, 8'd125, 8'd144, 8'd171, 8'd77, 8'd98, 8'd142, 8'd79, 8'd90, 8'd70, 8'd119, 8'd146, 8'd95, 8'd139, 8'd137, 8'd174, 8'd168, 8'd86, 8'd140, 8'd100, 8'd149, 8'd104, 8'd109, 8'd166, 8'd102, 8'd124, 8'd101, 8'd177, 8'd143, 8'd174, 8'd166, 8'd114, 8'd123, 8'd87, 8'd117, 8'd134, 8'd104, 8'd143, 8'd145, 8'd93, 8'd76, 8'd87, 8'd129, 8'd92, 8'd120, 8'd132, 8'd85, 8'd147, 8'd91, 8'd108, 8'd182, 8'd179, 8'd97, 8'd107, 8'd175, 8'd139, 8'd161, 8'd84, 8'd149, 8'd131, 8'd116, 8'd132, 8'd100, 8'd154, 8'd125, 8'd96, 8'd80, 8'd43, 8'd109, 8'd50, 8'd54, 8'd137, 8'd138, 8'd146, 8'd77, 8'd127, 8'd132, 8'd139, 8'd142, 8'd160, 8'd188, 8'd185, 8'd138, 8'd113, 8'd146, 8'd132, 8'd84, 8'd135, 8'd142, 8'd168, 8'd167, 8'd97, 8'd98, 8'd148, 8'd116, 8'd115, 8'd140, 8'd69, 8'd113, 8'd138, 8'd125, 8'd171, 8'd130, 8'd181, 8'd142, 8'd114, 8'd123, 8'd167, 8'd174, 8'd114, 8'd100, 8'd167, 8'd171, 8'd99, 8'd127, 8'd132, 8'd125, 8'd123, 8'd134, 8'd127, 8'd134, 8'd77, 8'd141, 8'd153, 8'd173, 8'd146, 8'd167, 8'd98, 8'd84, 8'd120, 8'd170, 8'd111, 8'd145, 8'd132, 8'd192, 8'd199, 8'd176, 8'd199, 8'd180, 8'd173, 8'd189, 8'd153, 8'd105, 8'd115, 8'd96, 8'd112, 8'd105, 8'd74, 8'd137, 8'd131, 8'd98, 8'd152, 8'd109, 8'd153, 8'd152, 8'd114, 8'd127, 8'd186, 8'd179, 8'd142, 8'd146, 8'd121, 8'd153, 8'd178, 8'd133, 8'd186, 8'd178, 8'd148, 8'd129, 8'd180, 8'd167, 8'd167, 8'd136, 8'd99, 8'd87, 8'd82, 8'd104, 8'd88, 8'd144, 8'd140, 8'd110, 8'd120, 8'd162, 8'd149, 8'd130, 8'd124, 8'd78, 8'd116, 8'd157, 8'd167, 8'd141, 8'd150, 8'd162, 8'd156, 8'd112, 8'd87, 8'd102, 8'd125, 8'd138, 8'd129, 8'd77, 8'd104, 8'd87, 8'd156})
) cell_0_94 (
    .clk(clk),
    .input_index(index_0_93_94),
    .input_value(value_0_93_94),
    .input_result(result_0_93_94),
    .input_enable(enable_0_93_94),
    .output_index(index_0_94_95),
    .output_value(value_0_94_95),
    .output_result(result_0_94_95),
    .output_enable(enable_0_94_95)
);

wire [10-1:0] index_0_95_96;
wire [`DATA_WIDTH-1:0] value_0_95_96;
wire [`DATA_WIDTH*4:0] result_0_95_96;
wire enable_0_95_96;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd169, 8'd153, 8'd98, 8'd99, 8'd59, 8'd65, 8'd90, 8'd68, 8'd97, 8'd74, 8'd57, 8'd146, 8'd101, 8'd132, 8'd111, 8'd114, 8'd122, 8'd153, 8'd156, 8'd145, 8'd69, 8'd73, 8'd98, 8'd134, 8'd117, 8'd96, 8'd113, 8'd72, 8'd167, 8'd102, 8'd67, 8'd169, 8'd149, 8'd125, 8'd118, 8'd98, 8'd63, 8'd93, 8'd80, 8'd135, 8'd117, 8'd154, 8'd125, 8'd134, 8'd123, 8'd73, 8'd122, 8'd158, 8'd76, 8'd166, 8'd125, 8'd174, 8'd98, 8'd165, 8'd165, 8'd116, 8'd150, 8'd137, 8'd147, 8'd160, 8'd191, 8'd155, 8'd124, 8'd135, 8'd88, 8'd145, 8'd113, 8'd172, 8'd84, 8'd105, 8'd80, 8'd58, 8'd73, 8'd138, 8'd123, 8'd48, 8'd127, 8'd85, 8'd62, 8'd95, 8'd123, 8'd163, 8'd155, 8'd133, 8'd113, 8'd110, 8'd150, 8'd92, 8'd136, 8'd178, 8'd162, 8'd173, 8'd100, 8'd180, 8'd94, 8'd91, 8'd106, 8'd76, 8'd132, 8'd72, 8'd82, 8'd76, 8'd63, 8'd108, 8'd51, 8'd47, 8'd122, 8'd83, 8'd70, 8'd99, 8'd144, 8'd159, 8'd75, 8'd141, 8'd152, 8'd141, 8'd179, 8'd184, 8'd147, 8'd90, 8'd155, 8'd116, 8'd166, 8'd104, 8'd164, 8'd156, 8'd157, 8'd75, 8'd125, 8'd95, 8'd106, 8'd142, 8'd83, 8'd89, 8'd135, 8'd95, 8'd114, 8'd72, 8'd93, 8'd164, 8'd84, 8'd143, 8'd127, 8'd118, 8'd139, 8'd124, 8'd109, 8'd145, 8'd100, 8'd128, 8'd156, 8'd88, 8'd104, 8'd95, 8'd107, 8'd109, 8'd90, 8'd95, 8'd77, 8'd64, 8'd73, 8'd64, 8'd105, 8'd124, 8'd141, 8'd51, 8'd107, 8'd125, 8'd128, 8'd87, 8'd149, 8'd138, 8'd136, 8'd165, 8'd181, 8'd124, 8'd94, 8'd93, 8'd94, 8'd73, 8'd99, 8'd147, 8'd163, 8'd133, 8'd156, 8'd154, 8'd163, 8'd128, 8'd150, 8'd104, 8'd99, 8'd119, 8'd97, 8'd138, 8'd152, 8'd88, 8'd97, 8'd145, 8'd155, 8'd93, 8'd172, 8'd89, 8'd73, 8'd73, 8'd78, 8'd76, 8'd123, 8'd109, 8'd147, 8'd112, 8'd78, 8'd116, 8'd159, 8'd68, 8'd124, 8'd90, 8'd93, 8'd123, 8'd95, 8'd132, 8'd93, 8'd101, 8'd154, 8'd71, 8'd132, 8'd54, 8'd98, 8'd141, 8'd161, 8'd127, 8'd122, 8'd158, 8'd158, 8'd81, 8'd131, 8'd159, 8'd103, 8'd113, 8'd88, 8'd119, 8'd82, 8'd153, 8'd116, 8'd142, 8'd80, 8'd109, 8'd87, 8'd130, 8'd122, 8'd138, 8'd72, 8'd68, 8'd136, 8'd79, 8'd83, 8'd158, 8'd134, 8'd68, 8'd59, 8'd151, 8'd133, 8'd132, 8'd119, 8'd156, 8'd81, 8'd175, 8'd123, 8'd95, 8'd133, 8'd90, 8'd178, 8'd124, 8'd129, 8'd152, 8'd79, 8'd103, 8'd59, 8'd63, 8'd72, 8'd125, 8'd141, 8'd104, 8'd72, 8'd65, 8'd111, 8'd123, 8'd61, 8'd107, 8'd85, 8'd99, 8'd74, 8'd162, 8'd114, 8'd106, 8'd148, 8'd156, 8'd134, 8'd77, 8'd87, 8'd70, 8'd107, 8'd103, 8'd110, 8'd102, 8'd115, 8'd44, 8'd133, 8'd78, 8'd114, 8'd60, 8'd88, 8'd60, 8'd87, 8'd94, 8'd86, 8'd123, 8'd97, 8'd149, 8'd65, 8'd82, 8'd116, 8'd138, 8'd113, 8'd126, 8'd135, 8'd88, 8'd144, 8'd93, 8'd71, 8'd78, 8'd65, 8'd128, 8'd125, 8'd54, 8'd118, 8'd65, 8'd83, 8'd59, 8'd34, 8'd142, 8'd104, 8'd75, 8'd101, 8'd127, 8'd110, 8'd150, 8'd114, 8'd83, 8'd121, 8'd79, 8'd153, 8'd113, 8'd142, 8'd107, 8'd126, 8'd142, 8'd111, 8'd119, 8'd102, 8'd109, 8'd122, 8'd146, 8'd158, 8'd169, 8'd94, 8'd118, 8'd37, 8'd129, 8'd111, 8'd65, 8'd115, 8'd138, 8'd71, 8'd141, 8'd73, 8'd96, 8'd164, 8'd73, 8'd113, 8'd167, 8'd141, 8'd103, 8'd124, 8'd156, 8'd114, 8'd169, 8'd104, 8'd153, 8'd80, 8'd65, 8'd83, 8'd157, 8'd74, 8'd88, 8'd119, 8'd99, 8'd87, 8'd156, 8'd128, 8'd133, 8'd92, 8'd143, 8'd85, 8'd118, 8'd102, 8'd150, 8'd170, 8'd124, 8'd199, 8'd116, 8'd137, 8'd165, 8'd160, 8'd118, 8'd164, 8'd160, 8'd114, 8'd83, 8'd91, 8'd66, 8'd120, 8'd174, 8'd91, 8'd77, 8'd82, 8'd99, 8'd135, 8'd153, 8'd119, 8'd104, 8'd59, 8'd80, 8'd126, 8'd165, 8'd100, 8'd136, 8'd122, 8'd169, 8'd161, 8'd139, 8'd156, 8'd184, 8'd140, 8'd161, 8'd116, 8'd53, 8'd110, 8'd132, 8'd112, 8'd156, 8'd159, 8'd152, 8'd104, 8'd108, 8'd64, 8'd109, 8'd77, 8'd34, 8'd134, 8'd101, 8'd73, 8'd149, 8'd124, 8'd134, 8'd197, 8'd149, 8'd142, 8'd121, 8'd181, 8'd150, 8'd92, 8'd124, 8'd64, 8'd38, 8'd55, 8'd139, 8'd157, 8'd122, 8'd175, 8'd185, 8'd146, 8'd132, 8'd95, 8'd119, 8'd71, 8'd122, 8'd119, 8'd123, 8'd47, 8'd149, 8'd123, 8'd155, 8'd130, 8'd176, 8'd141, 8'd153, 8'd156, 8'd97, 8'd83, 8'd116, 8'd38, 8'd100, 8'd146, 8'd154, 8'd94, 8'd175, 8'd227, 8'd211, 8'd177, 8'd164, 8'd154, 8'd153, 8'd91, 8'd137, 8'd107, 8'd87, 8'd33, 8'd128, 8'd157, 8'd151, 8'd189, 8'd131, 8'd160, 8'd136, 8'd81, 8'd59, 8'd96, 8'd106, 8'd121, 8'd59, 8'd128, 8'd155, 8'd85, 8'd165, 8'd170, 8'd184, 8'd185, 8'd140, 8'd148, 8'd163, 8'd122, 8'd68, 8'd108, 8'd70, 8'd120, 8'd102, 8'd113, 8'd110, 8'd106, 8'd160, 8'd92, 8'd120, 8'd145, 8'd87, 8'd57, 8'd39, 8'd97, 8'd56, 8'd96, 8'd122, 8'd125, 8'd167, 8'd126, 8'd208, 8'd187, 8'd116, 8'd165, 8'd158, 8'd107, 8'd161, 8'd85, 8'd145, 8'd100, 8'd68, 8'd147, 8'd140, 8'd75, 8'd152, 8'd153, 8'd123, 8'd95, 8'd69, 8'd106, 8'd82, 8'd101, 8'd95, 8'd152, 8'd132, 8'd108, 8'd96, 8'd193, 8'd192, 8'd143, 8'd101, 8'd112, 8'd177, 8'd150, 8'd113, 8'd161, 8'd90, 8'd91, 8'd117, 8'd109, 8'd99, 8'd149, 8'd120, 8'd140, 8'd147, 8'd88, 8'd46, 8'd74, 8'd107, 8'd88, 8'd142, 8'd117, 8'd150, 8'd74, 8'd188, 8'd161, 8'd102, 8'd174, 8'd144, 8'd154, 8'd96, 8'd180, 8'd168, 8'd133, 8'd81, 8'd159, 8'd81, 8'd126, 8'd155, 8'd115, 8'd63, 8'd80, 8'd71, 8'd136, 8'd97, 8'd85, 8'd43, 8'd85, 8'd143, 8'd125, 8'd147, 8'd145, 8'd123, 8'd143, 8'd168, 8'd89, 8'd123, 8'd171, 8'd86, 8'd127, 8'd87, 8'd99, 8'd95, 8'd159, 8'd68, 8'd113, 8'd133, 8'd102, 8'd121, 8'd59, 8'd54, 8'd119, 8'd116, 8'd87, 8'd62, 8'd80, 8'd128, 8'd120, 8'd160, 8'd106, 8'd128, 8'd137, 8'd155, 8'd141, 8'd77, 8'd174, 8'd164, 8'd82, 8'd66, 8'd93, 8'd67, 8'd124, 8'd87, 8'd105, 8'd37, 8'd72, 8'd112, 8'd108, 8'd48, 8'd95, 8'd90, 8'd136, 8'd143, 8'd121, 8'd113, 8'd157, 8'd96, 8'd158, 8'd72, 8'd108, 8'd139, 8'd133, 8'd68, 8'd80, 8'd75, 8'd116, 8'd90, 8'd48, 8'd47, 8'd84, 8'd36, 8'd11, 8'd80, 8'd67, 8'd56, 8'd60, 8'd121, 8'd122, 8'd63, 8'd73, 8'd94, 8'd90, 8'd141, 8'd131, 8'd97, 8'd132, 8'd106, 8'd131, 8'd113, 8'd130, 8'd66, 8'd125, 8'd61, 8'd76, 8'd126, 8'd123, 8'd112, 8'd52, 8'd87, 8'd59, 8'd84, 8'd89, 8'd51, 8'd83, 8'd95, 8'd109, 8'd131, 8'd68, 8'd144, 8'd93, 8'd159, 8'd105, 8'd170, 8'd165, 8'd106, 8'd97, 8'd143, 8'd96, 8'd120, 8'd72, 8'd111, 8'd98, 8'd162, 8'd124, 8'd88, 8'd125, 8'd168, 8'd80, 8'd127, 8'd101, 8'd102, 8'd112, 8'd112, 8'd156, 8'd124, 8'd84, 8'd94, 8'd167, 8'd106, 8'd85, 8'd140})
) cell_0_95 (
    .clk(clk),
    .input_index(index_0_94_95),
    .input_value(value_0_94_95),
    .input_result(result_0_94_95),
    .input_enable(enable_0_94_95),
    .output_index(index_0_95_96),
    .output_value(value_0_95_96),
    .output_result(result_0_95_96),
    .output_enable(enable_0_95_96)
);

wire [10-1:0] index_0_96_97;
wire [`DATA_WIDTH-1:0] value_0_96_97;
wire [`DATA_WIDTH*4:0] result_0_96_97;
wire enable_0_96_97;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd109, 8'd133, 8'd161, 8'd170, 8'd122, 8'd153, 8'd66, 8'd81, 8'd49, 8'd64, 8'd63, 8'd44, 8'd57, 8'd69, 8'd80, 8'd133, 8'd143, 8'd88, 8'd134, 8'd90, 8'd99, 8'd88, 8'd71, 8'd75, 8'd115, 8'd96, 8'd128, 8'd163, 8'd76, 8'd118, 8'd146, 8'd88, 8'd139, 8'd73, 8'd142, 8'd83, 8'd147, 8'd68, 8'd112, 8'd136, 8'd145, 8'd79, 8'd119, 8'd70, 8'd84, 8'd65, 8'd88, 8'd78, 8'd104, 8'd174, 8'd118, 8'd105, 8'd130, 8'd85, 8'd150, 8'd162, 8'd139, 8'd102, 8'd111, 8'd178, 8'd166, 8'd187, 8'd132, 8'd176, 8'd113, 8'd170, 8'd88, 8'd105, 8'd114, 8'd131, 8'd153, 8'd100, 8'd102, 8'd109, 8'd115, 8'd144, 8'd167, 8'd140, 8'd143, 8'd95, 8'd154, 8'd129, 8'd132, 8'd116, 8'd138, 8'd71, 8'd92, 8'd65, 8'd139, 8'd125, 8'd115, 8'd121, 8'd172, 8'd148, 8'd150, 8'd94, 8'd158, 8'd119, 8'd174, 8'd108, 8'd153, 8'd199, 8'd105, 8'd119, 8'd128, 8'd108, 8'd170, 8'd176, 8'd130, 8'd98, 8'd145, 8'd144, 8'd111, 8'd83, 8'd80, 8'd145, 8'd142, 8'd90, 8'd109, 8'd135, 8'd132, 8'd113, 8'd86, 8'd90, 8'd111, 8'd94, 8'd135, 8'd116, 8'd143, 8'd84, 8'd153, 8'd94, 8'd106, 8'd125, 8'd158, 8'd150, 8'd127, 8'd100, 8'd170, 8'd129, 8'd154, 8'd131, 8'd124, 8'd90, 8'd77, 8'd112, 8'd77, 8'd155, 8'd87, 8'd109, 8'd97, 8'd141, 8'd143, 8'd109, 8'd105, 8'd153, 8'd136, 8'd110, 8'd98, 8'd122, 8'd106, 8'd71, 8'd150, 8'd147, 8'd152, 8'd112, 8'd97, 8'd89, 8'd91, 8'd152, 8'd57, 8'd112, 8'd123, 8'd117, 8'd122, 8'd115, 8'd145, 8'd110, 8'd83, 8'd115, 8'd104, 8'd111, 8'd129, 8'd79, 8'd147, 8'd97, 8'd108, 8'd66, 8'd75, 8'd129, 8'd93, 8'd85, 8'd99, 8'd152, 8'd168, 8'd110, 8'd169, 8'd55, 8'd102, 8'd123, 8'd103, 8'd147, 8'd72, 8'd162, 8'd98, 8'd112, 8'd114, 8'd168, 8'd102, 8'd161, 8'd102, 8'd105, 8'd148, 8'd90, 8'd91, 8'd151, 8'd98, 8'd71, 8'd81, 8'd79, 8'd171, 8'd88, 8'd157, 8'd163, 8'd79, 8'd70, 8'd107, 8'd120, 8'd114, 8'd75, 8'd153, 8'd153, 8'd178, 8'd93, 8'd89, 8'd172, 8'd145, 8'd154, 8'd98, 8'd114, 8'd88, 8'd124, 8'd126, 8'd101, 8'd69, 8'd139, 8'd71, 8'd82, 8'd187, 8'd132, 8'd79, 8'd92, 8'd62, 8'd134, 8'd36, 8'd81, 8'd125, 8'd108, 8'd112, 8'd144, 8'd120, 8'd181, 8'd118, 8'd139, 8'd134, 8'd81, 8'd108, 8'd81, 8'd82, 8'd78, 8'd155, 8'd148, 8'd77, 8'd101, 8'd81, 8'd160, 8'd140, 8'd147, 8'd93, 8'd155, 8'd117, 8'd121, 8'd99, 8'd120, 8'd103, 8'd96, 8'd118, 8'd149, 8'd87, 8'd137, 8'd124, 8'd138, 8'd112, 8'd86, 8'd101, 8'd82, 8'd86, 8'd88, 8'd135, 8'd88, 8'd61, 8'd69, 8'd142, 8'd80, 8'd120, 8'd110, 8'd101, 8'd75, 8'd127, 8'd84, 8'd46, 8'd131, 8'd81, 8'd132, 8'd115, 8'd105, 8'd125, 8'd154, 8'd112, 8'd166, 8'd138, 8'd152, 8'd76, 8'd122, 8'd148, 8'd152, 8'd144, 8'd124, 8'd66, 8'd134, 8'd77, 8'd123, 8'd135, 8'd77, 8'd81, 8'd82, 8'd135, 8'd41, 8'd125, 8'd129, 8'd152, 8'd161, 8'd136, 8'd144, 8'd135, 8'd96, 8'd111, 8'd95, 8'd96, 8'd131, 8'd86, 8'd111, 8'd200, 8'd197, 8'd181, 8'd164, 8'd158, 8'd139, 8'd109, 8'd138, 8'd133, 8'd112, 8'd98, 8'd96, 8'd112, 8'd49, 8'd74, 8'd126, 8'd152, 8'd134, 8'd168, 8'd166, 8'd160, 8'd138, 8'd113, 8'd103, 8'd163, 8'd108, 8'd153, 8'd152, 8'd197, 8'd172, 8'd189, 8'd95, 8'd179, 8'd132, 8'd128, 8'd142, 8'd121, 8'd127, 8'd127, 8'd101, 8'd118, 8'd45, 8'd51, 8'd40, 8'd87, 8'd103, 8'd79, 8'd139, 8'd127, 8'd91, 8'd170, 8'd134, 8'd126, 8'd150, 8'd129, 8'd188, 8'd208, 8'd125, 8'd103, 8'd154, 8'd189, 8'd203, 8'd178, 8'd134, 8'd121, 8'd60, 8'd153, 8'd140, 8'd130, 8'd85, 8'd135, 8'd69, 8'd79, 8'd81, 8'd118, 8'd148, 8'd133, 8'd122, 8'd151, 8'd141, 8'd118, 8'd198, 8'd182, 8'd166, 8'd216, 8'd201, 8'd150, 8'd110, 8'd171, 8'd216, 8'd159, 8'd89, 8'd110, 8'd122, 8'd119, 8'd81, 8'd88, 8'd114, 8'd124, 8'd146, 8'd129, 8'd83, 8'd119, 8'd79, 8'd121, 8'd148, 8'd149, 8'd132, 8'd150, 8'd92, 8'd160, 8'd167, 8'd175, 8'd175, 8'd128, 8'd110, 8'd186, 8'd151, 8'd168, 8'd139, 8'd105, 8'd59, 8'd76, 8'd161, 8'd143, 8'd193, 8'd170, 8'd205, 8'd113, 8'd128, 8'd114, 8'd62, 8'd65, 8'd115, 8'd47, 8'd77, 8'd56, 8'd84, 8'd99, 8'd146, 8'd164, 8'd77, 8'd167, 8'd119, 8'd146, 8'd126, 8'd92, 8'd138, 8'd114, 8'd88, 8'd148, 8'd81, 8'd73, 8'd125, 8'd219, 8'd205, 8'd86, 8'd163, 8'd154, 8'd136, 8'd143, 8'd82, 8'd108, 8'd51, 8'd47, 8'd79, 8'd102, 8'd161, 8'd137, 8'd74, 8'd61, 8'd161, 8'd106, 8'd152, 8'd70, 8'd85, 8'd45, 8'd96, 8'd77, 8'd74, 8'd104, 8'd136, 8'd124, 8'd190, 8'd91, 8'd85, 8'd103, 8'd113, 8'd151, 8'd90, 8'd98, 8'd127, 8'd134, 8'd109, 8'd106, 8'd105, 8'd157, 8'd81, 8'd106, 8'd110, 8'd76, 8'd77, 8'd85, 8'd34, 8'd97, 8'd60, 8'd92, 8'd113, 8'd165, 8'd142, 8'd108, 8'd189, 8'd109, 8'd146, 8'd98, 8'd73, 8'd151, 8'd107, 8'd96, 8'd89, 8'd83, 8'd156, 8'd82, 8'd97, 8'd102, 8'd145, 8'd124, 8'd119, 8'd143, 8'd125, 8'd64, 8'd121, 8'd138, 8'd147, 8'd130, 8'd144, 8'd95, 8'd127, 8'd163, 8'd152, 8'd147, 8'd132, 8'd122, 8'd111, 8'd104, 8'd124, 8'd145, 8'd116, 8'd145, 8'd120, 8'd107, 8'd93, 8'd72, 8'd119, 8'd151, 8'd129, 8'd147, 8'd61, 8'd84, 8'd79, 8'd140, 8'd113, 8'd120, 8'd104, 8'd104, 8'd186, 8'd194, 8'd197, 8'd103, 8'd151, 8'd81, 8'd150, 8'd168, 8'd105, 8'd76, 8'd138, 8'd139, 8'd85, 8'd63, 8'd62, 8'd127, 8'd103, 8'd139, 8'd87, 8'd147, 8'd163, 8'd99, 8'd97, 8'd102, 8'd150, 8'd139, 8'd112, 8'd162, 8'd113, 8'd93, 8'd164, 8'd158, 8'd138, 8'd125, 8'd141, 8'd175, 8'd104, 8'd87, 8'd153, 8'd152, 8'd133, 8'd92, 8'd86, 8'd113, 8'd103, 8'd150, 8'd150, 8'd142, 8'd115, 8'd109, 8'd84, 8'd90, 8'd144, 8'd114, 8'd121, 8'd73, 8'd170, 8'd164, 8'd100, 8'd99, 8'd144, 8'd128, 8'd179, 8'd179, 8'd140, 8'd94, 8'd146, 8'd112, 8'd112, 8'd61, 8'd82, 8'd97, 8'd148, 8'd81, 8'd77, 8'd120, 8'd166, 8'd159, 8'd176, 8'd102, 8'd148, 8'd143, 8'd82, 8'd148, 8'd124, 8'd66, 8'd144, 8'd163, 8'd177, 8'd138, 8'd120, 8'd136, 8'd161, 8'd78, 8'd149, 8'd81, 8'd109, 8'd122, 8'd160, 8'd166, 8'd156, 8'd109, 8'd133, 8'd96, 8'd98, 8'd84, 8'd137, 8'd70, 8'd131, 8'd101, 8'd162, 8'd97, 8'd86, 8'd132, 8'd134, 8'd91, 8'd88, 8'd150, 8'd139, 8'd94, 8'd168, 8'd118, 8'd66, 8'd79, 8'd97, 8'd111, 8'd178, 8'd138, 8'd166, 8'd167, 8'd76, 8'd92, 8'd79, 8'd150, 8'd100, 8'd113, 8'd102, 8'd123, 8'd156, 8'd78, 8'd99, 8'd106, 8'd152, 8'd101, 8'd72, 8'd152, 8'd143, 8'd102, 8'd145, 8'd108, 8'd162, 8'd127, 8'd92, 8'd132, 8'd91, 8'd134, 8'd140, 8'd120, 8'd123, 8'd95, 8'd144, 8'd165, 8'd91, 8'd98, 8'd88, 8'd109, 8'd85})
) cell_0_96 (
    .clk(clk),
    .input_index(index_0_95_96),
    .input_value(value_0_95_96),
    .input_result(result_0_95_96),
    .input_enable(enable_0_95_96),
    .output_index(index_0_96_97),
    .output_value(value_0_96_97),
    .output_result(result_0_96_97),
    .output_enable(enable_0_96_97)
);

wire [10-1:0] index_0_97_98;
wire [`DATA_WIDTH-1:0] value_0_97_98;
wire [`DATA_WIDTH*4:0] result_0_97_98;
wire enable_0_97_98;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd91, 8'd105, 8'd120, 8'd164, 8'd84, 8'd86, 8'd146, 8'd104, 8'd101, 8'd145, 8'd47, 8'd148, 8'd72, 8'd133, 8'd51, 8'd119, 8'd133, 8'd77, 8'd102, 8'd93, 8'd82, 8'd113, 8'd159, 8'd123, 8'd115, 8'd82, 8'd124, 8'd146, 8'd167, 8'd111, 8'd67, 8'd90, 8'd104, 8'd70, 8'd158, 8'd117, 8'd163, 8'd182, 8'd130, 8'd83, 8'd98, 8'd120, 8'd179, 8'd137, 8'd133, 8'd131, 8'd156, 8'd120, 8'd149, 8'd138, 8'd126, 8'd175, 8'd112, 8'd153, 8'd132, 8'd131, 8'd75, 8'd66, 8'd130, 8'd152, 8'd100, 8'd179, 8'd195, 8'd115, 8'd97, 8'd90, 8'd177, 8'd176, 8'd82, 8'd96, 8'd170, 8'd121, 8'd177, 8'd122, 8'd189, 8'd104, 8'd171, 8'd177, 8'd168, 8'd153, 8'd74, 8'd88, 8'd83, 8'd107, 8'd110, 8'd121, 8'd86, 8'd90, 8'd167, 8'd91, 8'd145, 8'd99, 8'd99, 8'd86, 8'd75, 8'd113, 8'd65, 8'd88, 8'd154, 8'd154, 8'd85, 8'd133, 8'd134, 8'd139, 8'd98, 8'd94, 8'd168, 8'd84, 8'd128, 8'd167, 8'd116, 8'd137, 8'd77, 8'd144, 8'd107, 8'd128, 8'd162, 8'd148, 8'd102, 8'd165, 8'd84, 8'd107, 8'd112, 8'd126, 8'd145, 8'd90, 8'd113, 8'd82, 8'd116, 8'd101, 8'd92, 8'd138, 8'd142, 8'd59, 8'd87, 8'd65, 8'd130, 8'd135, 8'd159, 8'd126, 8'd113, 8'd90, 8'd140, 8'd146, 8'd144, 8'd156, 8'd92, 8'd78, 8'd142, 8'd129, 8'd139, 8'd102, 8'd75, 8'd156, 8'd130, 8'd150, 8'd144, 8'd75, 8'd91, 8'd64, 8'd55, 8'd89, 8'd70, 8'd62, 8'd135, 8'd134, 8'd140, 8'd78, 8'd111, 8'd122, 8'd148, 8'd68, 8'd147, 8'd147, 8'd151, 8'd148, 8'd103, 8'd85, 8'd99, 8'd85, 8'd151, 8'd169, 8'd115, 8'd64, 8'd102, 8'd114, 8'd130, 8'd138, 8'd86, 8'd150, 8'd81, 8'd68, 8'd78, 8'd68, 8'd131, 8'd83, 8'd88, 8'd121, 8'd81, 8'd141, 8'd117, 8'd150, 8'd151, 8'd137, 8'd149, 8'd109, 8'd160, 8'd119, 8'd72, 8'd66, 8'd142, 8'd161, 8'd113, 8'd100, 8'd142, 8'd57, 8'd132, 8'd71, 8'd142, 8'd63, 8'd119, 8'd96, 8'd112, 8'd75, 8'd121, 8'd124, 8'd114, 8'd140, 8'd130, 8'd84, 8'd104, 8'd159, 8'd109, 8'd99, 8'd115, 8'd151, 8'd129, 8'd140, 8'd68, 8'd123, 8'd62, 8'd132, 8'd137, 8'd140, 8'd140, 8'd70, 8'd84, 8'd67, 8'd142, 8'd158, 8'd154, 8'd83, 8'd78, 8'd135, 8'd121, 8'd126, 8'd80, 8'd149, 8'd106, 8'd74, 8'd99, 8'd85, 8'd170, 8'd115, 8'd157, 8'd151, 8'd152, 8'd108, 8'd136, 8'd114, 8'd82, 8'd62, 8'd137, 8'd112, 8'd49, 8'd57, 8'd129, 8'd122, 8'd127, 8'd125, 8'd133, 8'd87, 8'd99, 8'd127, 8'd99, 8'd153, 8'd79, 8'd121, 8'd82, 8'd105, 8'd87, 8'd152, 8'd136, 8'd128, 8'd149, 8'd143, 8'd160, 8'd82, 8'd86, 8'd102, 8'd115, 8'd103, 8'd101, 8'd72, 8'd147, 8'd113, 8'd152, 8'd109, 8'd146, 8'd42, 8'd71, 8'd123, 8'd71, 8'd109, 8'd114, 8'd114, 8'd163, 8'd158, 8'd134, 8'd142, 8'd112, 8'd117, 8'd148, 8'd143, 8'd106, 8'd94, 8'd107, 8'd168, 8'd140, 8'd125, 8'd138, 8'd107, 8'd83, 8'd137, 8'd141, 8'd128, 8'd75, 8'd77, 8'd81, 8'd105, 8'd159, 8'd118, 8'd167, 8'd78, 8'd73, 8'd166, 8'd132, 8'd161, 8'd169, 8'd145, 8'd140, 8'd154, 8'd109, 8'd99, 8'd90, 8'd118, 8'd101, 8'd87, 8'd64, 8'd143, 8'd137, 8'd156, 8'd169, 8'd80, 8'd149, 8'd48, 8'd114, 8'd98, 8'd116, 8'd89, 8'd119, 8'd120, 8'd79, 8'd169, 8'd93, 8'd105, 8'd158, 8'd124, 8'd181, 8'd120, 8'd134, 8'd170, 8'd125, 8'd169, 8'd118, 8'd119, 8'd119, 8'd154, 8'd152, 8'd76, 8'd112, 8'd142, 8'd117, 8'd63, 8'd75, 8'd135, 8'd171, 8'd136, 8'd105, 8'd108, 8'd134, 8'd85, 8'd107, 8'd152, 8'd149, 8'd166, 8'd214, 8'd143, 8'd142, 8'd99, 8'd129, 8'd92, 8'd159, 8'd167, 8'd110, 8'd167, 8'd128, 8'd143, 8'd110, 8'd157, 8'd128, 8'd52, 8'd126, 8'd73, 8'd119, 8'd158, 8'd136, 8'd91, 8'd124, 8'd136, 8'd121, 8'd171, 8'd144, 8'd140, 8'd214, 8'd216, 8'd151, 8'd164, 8'd190, 8'd193, 8'd107, 8'd142, 8'd192, 8'd78, 8'd102, 8'd75, 8'd69, 8'd138, 8'd87, 8'd165, 8'd133, 8'd155, 8'd138, 8'd106, 8'd124, 8'd109, 8'd132, 8'd121, 8'd134, 8'd84, 8'd148, 8'd118, 8'd168, 8'd197, 8'd121, 8'd186, 8'd168, 8'd113, 8'd152, 8'd141, 8'd106, 8'd94, 8'd44, 8'd50, 8'd55, 8'd145, 8'd140, 8'd106, 8'd161, 8'd130, 8'd117, 8'd65, 8'd66, 8'd110, 8'd92, 8'd124, 8'd89, 8'd44, 8'd82, 8'd147, 8'd161, 8'd103, 8'd127, 8'd89, 8'd86, 8'd102, 8'd154, 8'd107, 8'd61, 8'd100, 8'd127, 8'd86, 8'd87, 8'd107, 8'd109, 8'd123, 8'd191, 8'd180, 8'd91, 8'd77, 8'd126, 8'd87, 8'd105, 8'd46, 8'd43, 8'd90, 8'd79, 8'd122, 8'd150, 8'd115, 8'd139, 8'd69, 8'd158, 8'd93, 8'd147, 8'd63, 8'd75, 8'd94, 8'd42, 8'd58, 8'd74, 8'd140, 8'd105, 8'd180, 8'd111, 8'd147, 8'd73, 8'd53, 8'd85, 8'd112, 8'd108, 8'd147, 8'd129, 8'd77, 8'd101, 8'd112, 8'd86, 8'd124, 8'd123, 8'd101, 8'd91, 8'd126, 8'd67, 8'd63, 8'd118, 8'd57, 8'd66, 8'd81, 8'd134, 8'd80, 8'd96, 8'd171, 8'd121, 8'd94, 8'd148, 8'd62, 8'd134, 8'd136, 8'd61, 8'd114, 8'd88, 8'd174, 8'd128, 8'd116, 8'd160, 8'd142, 8'd83, 8'd93, 8'd84, 8'd132, 8'd90, 8'd99, 8'd59, 8'd97, 8'd75, 8'd80, 8'd95, 8'd71, 8'd96, 8'd106, 8'd173, 8'd124, 8'd141, 8'd101, 8'd150, 8'd114, 8'd106, 8'd73, 8'd132, 8'd82, 8'd165, 8'd159, 8'd87, 8'd87, 8'd74, 8'd55, 8'd64, 8'd88, 8'd145, 8'd45, 8'd85, 8'd101, 8'd92, 8'd83, 8'd137, 8'd165, 8'd124, 8'd136, 8'd168, 8'd166, 8'd139, 8'd131, 8'd147, 8'd92, 8'd122, 8'd125, 8'd91, 8'd124, 8'd56, 8'd106, 8'd150, 8'd151, 8'd118, 8'd145, 8'd64, 8'd106, 8'd87, 8'd69, 8'd92, 8'd97, 8'd89, 8'd121, 8'd71, 8'd123, 8'd161, 8'd157, 8'd179, 8'd210, 8'd146, 8'd206, 8'd198, 8'd189, 8'd129, 8'd167, 8'd111, 8'd153, 8'd143, 8'd148, 8'd123, 8'd120, 8'd126, 8'd90, 8'd101, 8'd110, 8'd70, 8'd70, 8'd94, 8'd86, 8'd70, 8'd145, 8'd95, 8'd168, 8'd126, 8'd168, 8'd124, 8'd152, 8'd192, 8'd184, 8'd160, 8'd187, 8'd169, 8'd145, 8'd84, 8'd147, 8'd154, 8'd122, 8'd66, 8'd136, 8'd78, 8'd100, 8'd154, 8'd112, 8'd159, 8'd169, 8'd141, 8'd87, 8'd148, 8'd93, 8'd106, 8'd160, 8'd73, 8'd169, 8'd154, 8'd80, 8'd100, 8'd159, 8'd185, 8'd155, 8'd182, 8'd181, 8'd135, 8'd82, 8'd164, 8'd176, 8'd159, 8'd125, 8'd139, 8'd128, 8'd108, 8'd120, 8'd123, 8'd154, 8'd125, 8'd172, 8'd99, 8'd139, 8'd112, 8'd99, 8'd129, 8'd83, 8'd149, 8'd163, 8'd115, 8'd102, 8'd150, 8'd163, 8'd158, 8'd136, 8'd81, 8'd99, 8'd75, 8'd142, 8'd150, 8'd127, 8'd115, 8'd161, 8'd138, 8'd138, 8'd99, 8'd163, 8'd148, 8'd126, 8'd138, 8'd120, 8'd156, 8'd121, 8'd124, 8'd92, 8'd120, 8'd132, 8'd130, 8'd90, 8'd75, 8'd90, 8'd118, 8'd152, 8'd109, 8'd102, 8'd111, 8'd99, 8'd154, 8'd135, 8'd158, 8'd146, 8'd102, 8'd103, 8'd81, 8'd119, 8'd124, 8'd166, 8'd156, 8'd83, 8'd138, 8'd130})
) cell_0_97 (
    .clk(clk),
    .input_index(index_0_96_97),
    .input_value(value_0_96_97),
    .input_result(result_0_96_97),
    .input_enable(enable_0_96_97),
    .output_index(index_0_97_98),
    .output_value(value_0_97_98),
    .output_result(result_0_97_98),
    .output_enable(enable_0_97_98)
);

wire [10-1:0] index_0_98_99;
wire [`DATA_WIDTH-1:0] value_0_98_99;
wire [`DATA_WIDTH*4:0] result_0_98_99;
wire enable_0_98_99;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd89, 8'd124, 8'd123, 8'd80, 8'd155, 8'd159, 8'd122, 8'd152, 8'd114, 8'd189, 8'd165, 8'd117, 8'd171, 8'd185, 8'd154, 8'd162, 8'd126, 8'd147, 8'd163, 8'd156, 8'd155, 8'd163, 8'd108, 8'd130, 8'd120, 8'd116, 8'd144, 8'd161, 8'd111, 8'd154, 8'd113, 8'd120, 8'd130, 8'd127, 8'd112, 8'd147, 8'd178, 8'd105, 8'd143, 8'd130, 8'd127, 8'd171, 8'd158, 8'd125, 8'd118, 8'd118, 8'd145, 8'd128, 8'd178, 8'd170, 8'd142, 8'd128, 8'd93, 8'd152, 8'd167, 8'd109, 8'd132, 8'd111, 8'd131, 8'd121, 8'd131, 8'd133, 8'd102, 8'd121, 8'd104, 8'd110, 8'd163, 8'd168, 8'd99, 8'd95, 8'd115, 8'd115, 8'd92, 8'd119, 8'd100, 8'd96, 8'd172, 8'd116, 8'd86, 8'd124, 8'd171, 8'd79, 8'd101, 8'd139, 8'd70, 8'd111, 8'd123, 8'd143, 8'd114, 8'd73, 8'd150, 8'd125, 8'd98, 8'd71, 8'd166, 8'd115, 8'd111, 8'd138, 8'd95, 8'd168, 8'd87, 8'd72, 8'd138, 8'd94, 8'd163, 8'd168, 8'd131, 8'd110, 8'd79, 8'd159, 8'd157, 8'd71, 8'd72, 8'd86, 8'd91, 8'd66, 8'd65, 8'd85, 8'd74, 8'd140, 8'd110, 8'd72, 8'd144, 8'd101, 8'd160, 8'd97, 8'd144, 8'd105, 8'd66, 8'd134, 8'd98, 8'd102, 8'd149, 8'd129, 8'd113, 8'd88, 8'd59, 8'd109, 8'd89, 8'd70, 8'd133, 8'd118, 8'd66, 8'd53, 8'd90, 8'd89, 8'd108, 8'd114, 8'd82, 8'd112, 8'd68, 8'd140, 8'd176, 8'd111, 8'd148, 8'd149, 8'd58, 8'd141, 8'd128, 8'd132, 8'd90, 8'd107, 8'd130, 8'd39, 8'd29, 8'd60, 8'd99, 8'd71, 8'd129, 8'd148, 8'd96, 8'd89, 8'd71, 8'd104, 8'd97, 8'd95, 8'd84, 8'd140, 8'd74, 8'd142, 8'd146, 8'd143, 8'd146, 8'd100, 8'd92, 8'd130, 8'd96, 8'd134, 8'd142, 8'd114, 8'd54, 8'd48, 8'd31, 8'd106, 8'd157, 8'd111, 8'd156, 8'd143, 8'd81, 8'd128, 8'd57, 8'd107, 8'd135, 8'd94, 8'd85, 8'd98, 8'd118, 8'd69, 8'd76, 8'd136, 8'd184, 8'd153, 8'd166, 8'd74, 8'd94, 8'd95, 8'd76, 8'd94, 8'd48, 8'd102, 8'd55, 8'd130, 8'd75, 8'd91, 8'd87, 8'd64, 8'd64, 8'd51, 8'd112, 8'd94, 8'd126, 8'd115, 8'd123, 8'd74, 8'd117, 8'd147, 8'd87, 8'd168, 8'd85, 8'd140, 8'd123, 8'd145, 8'd121, 8'd54, 8'd122, 8'd66, 8'd77, 8'd45, 8'd71, 8'd123, 8'd129, 8'd74, 8'd135, 8'd87, 8'd77, 8'd90, 8'd126, 8'd54, 8'd109, 8'd104, 8'd68, 8'd74, 8'd96, 8'd122, 8'd155, 8'd96, 8'd171, 8'd147, 8'd154, 8'd176, 8'd137, 8'd123, 8'd78, 8'd70, 8'd71, 8'd21, 8'd46, 8'd69, 8'd146, 8'd90, 8'd135, 8'd133, 8'd127, 8'd143, 8'd93, 8'd93, 8'd75, 8'd139, 8'd91, 8'd75, 8'd116, 8'd114, 8'd105, 8'd123, 8'd113, 8'd164, 8'd139, 8'd96, 8'd183, 8'd84, 8'd150, 8'd59, 8'd86, 8'd106, 8'd109, 8'd80, 8'd161, 8'd85, 8'd145, 8'd103, 8'd92, 8'd109, 8'd157, 8'd143, 8'd158, 8'd136, 8'd94, 8'd96, 8'd168, 8'd164, 8'd159, 8'd135, 8'd119, 8'd116, 8'd153, 8'd172, 8'd109, 8'd97, 8'd113, 8'd149, 8'd126, 8'd96, 8'd135, 8'd72, 8'd153, 8'd163, 8'd94, 8'd49, 8'd81, 8'd155, 8'd86, 8'd146, 8'd115, 8'd130, 8'd105, 8'd180, 8'd96, 8'd137, 8'd96, 8'd155, 8'd83, 8'd128, 8'd111, 8'd153, 8'd138, 8'd135, 8'd133, 8'd83, 8'd92, 8'd127, 8'd94, 8'd92, 8'd103, 8'd110, 8'd130, 8'd78, 8'd123, 8'd142, 8'd117, 8'd127, 8'd95, 8'd95, 8'd110, 8'd177, 8'd105, 8'd100, 8'd115, 8'd123, 8'd80, 8'd76, 8'd100, 8'd159, 8'd130, 8'd169, 8'd163, 8'd201, 8'd190, 8'd165, 8'd175, 8'd155, 8'd115, 8'd100, 8'd151, 8'd94, 8'd78, 8'd118, 8'd172, 8'd154, 8'd162, 8'd180, 8'd159, 8'd142, 8'd117, 8'd99, 8'd128, 8'd69, 8'd72, 8'd112, 8'd142, 8'd155, 8'd135, 8'd188, 8'd192, 8'd198, 8'd169, 8'd140, 8'd133, 8'd126, 8'd119, 8'd147, 8'd110, 8'd112, 8'd103, 8'd133, 8'd140, 8'd157, 8'd128, 8'd91, 8'd85, 8'd104, 8'd143, 8'd139, 8'd62, 8'd102, 8'd60, 8'd183, 8'd114, 8'd184, 8'd126, 8'd144, 8'd208, 8'd207, 8'd141, 8'd95, 8'd97, 8'd169, 8'd152, 8'd122, 8'd148, 8'd52, 8'd86, 8'd122, 8'd151, 8'd198, 8'd119, 8'd169, 8'd125, 8'd143, 8'd159, 8'd121, 8'd85, 8'd135, 8'd188, 8'd156, 8'd145, 8'd176, 8'd165, 8'd215, 8'd209, 8'd98, 8'd96, 8'd156, 8'd135, 8'd126, 8'd128, 8'd96, 8'd93, 8'd43, 8'd23, 8'd69, 8'd138, 8'd137, 8'd119, 8'd92, 8'd106, 8'd135, 8'd84, 8'd161, 8'd123, 8'd64, 8'd91, 8'd132, 8'd179, 8'd201, 8'd169, 8'd152, 8'd107, 8'd100, 8'd100, 8'd119, 8'd113, 8'd107, 8'd120, 8'd130, 8'd77, 8'd147, 8'd115, 8'd128, 8'd155, 8'd92, 8'd98, 8'd146, 8'd138, 8'd86, 8'd94, 8'd57, 8'd124, 8'd92, 8'd130, 8'd93, 8'd188, 8'd160, 8'd93, 8'd114, 8'd180, 8'd138, 8'd103, 8'd141, 8'd120, 8'd169, 8'd134, 8'd88, 8'd92, 8'd156, 8'd137, 8'd142, 8'd126, 8'd134, 8'd173, 8'd91, 8'd159, 8'd104, 8'd71, 8'd149, 8'd136, 8'd140, 8'd140, 8'd143, 8'd128, 8'd117, 8'd136, 8'd114, 8'd132, 8'd108, 8'd76, 8'd129, 8'd122, 8'd117, 8'd82, 8'd145, 8'd151, 8'd148, 8'd92, 8'd120, 8'd150, 8'd116, 8'd85, 8'd110, 8'd116, 8'd94, 8'd107, 8'd59, 8'd122, 8'd102, 8'd112, 8'd158, 8'd165, 8'd145, 8'd175, 8'd81, 8'd94, 8'd156, 8'd118, 8'd134, 8'd143, 8'd125, 8'd93, 8'd120, 8'd113, 8'd121, 8'd137, 8'd152, 8'd119, 8'd131, 8'd163, 8'd110, 8'd157, 8'd64, 8'd78, 8'd145, 8'd68, 8'd117, 8'd67, 8'd69, 8'd158, 8'd91, 8'd97, 8'd151, 8'd94, 8'd101, 8'd148, 8'd130, 8'd154, 8'd169, 8'd78, 8'd143, 8'd96, 8'd95, 8'd182, 8'd203, 8'd143, 8'd128, 8'd114, 8'd106, 8'd91, 8'd97, 8'd103, 8'd134, 8'd55, 8'd147, 8'd142, 8'd85, 8'd80, 8'd110, 8'd144, 8'd74, 8'd78, 8'd133, 8'd91, 8'd128, 8'd102, 8'd78, 8'd80, 8'd133, 8'd84, 8'd138, 8'd108, 8'd198, 8'd192, 8'd192, 8'd205, 8'd168, 8'd157, 8'd154, 8'd88, 8'd70, 8'd96, 8'd62, 8'd88, 8'd122, 8'd74, 8'd50, 8'd72, 8'd114, 8'd93, 8'd145, 8'd73, 8'd135, 8'd135, 8'd85, 8'd158, 8'd110, 8'd163, 8'd168, 8'd173, 8'd94, 8'd186, 8'd134, 8'd180, 8'd147, 8'd109, 8'd173, 8'd111, 8'd138, 8'd156, 8'd78, 8'd143, 8'd101, 8'd115, 8'd77, 8'd106, 8'd150, 8'd105, 8'd100, 8'd86, 8'd149, 8'd152, 8'd164, 8'd108, 8'd158, 8'd160, 8'd75, 8'd67, 8'd168, 8'd173, 8'd149, 8'd165, 8'd185, 8'd186, 8'd111, 8'd105, 8'd162, 8'd120, 8'd85, 8'd99, 8'd162, 8'd156, 8'd176, 8'd160, 8'd129, 8'd132, 8'd109, 8'd132, 8'd134, 8'd70, 8'd154, 8'd126, 8'd153, 8'd78, 8'd109, 8'd132, 8'd117, 8'd117, 8'd84, 8'd147, 8'd119, 8'd102, 8'd164, 8'd167, 8'd136, 8'd116, 8'd133, 8'd151, 8'd163, 8'd167, 8'd131, 8'd152, 8'd162, 8'd137, 8'd114, 8'd126, 8'd88, 8'd142, 8'd138, 8'd149, 8'd131, 8'd127, 8'd83, 8'd148, 8'd85, 8'd106, 8'd166, 8'd81, 8'd71, 8'd102, 8'd162, 8'd141, 8'd70, 8'd75, 8'd116, 8'd168, 8'd100, 8'd132, 8'd111, 8'd110, 8'd134, 8'd136, 8'd156, 8'd139, 8'd136, 8'd124, 8'd138, 8'd128, 8'd121})
) cell_0_98 (
    .clk(clk),
    .input_index(index_0_97_98),
    .input_value(value_0_97_98),
    .input_result(result_0_97_98),
    .input_enable(enable_0_97_98),
    .output_index(index_0_98_99),
    .output_value(value_0_98_99),
    .output_result(result_0_98_99),
    .output_enable(enable_0_98_99)
);

wire [10-1:0] index_0_99_100;
wire [`DATA_WIDTH-1:0] value_0_99_100;
wire [`DATA_WIDTH*4:0] result_0_99_100;
wire enable_0_99_100;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(10),
    .WEIGHT_AMOUNT(784),
    .WEIGHT_OFFSET(120),
    .INPUT_OFFSET(0),
    .WEIGHTS({8'd133, 8'd122, 8'd98, 8'd150, 8'd134, 8'd99, 8'd134, 8'd104, 8'd126, 8'd129, 8'd145, 8'd141, 8'd95, 8'd171, 8'd208, 8'd165, 8'd169, 8'd123, 8'd151, 8'd98, 8'd90, 8'd109, 8'd178, 8'd96, 8'd140, 8'd81, 8'd101, 8'd123, 8'd78, 8'd133, 8'd113, 8'd157, 8'd165, 8'd122, 8'd146, 8'd140, 8'd119, 8'd187, 8'd116, 8'd106, 8'd163, 8'd175, 8'd89, 8'd133, 8'd157, 8'd88, 8'd96, 8'd115, 8'd133, 8'd86, 8'd150, 8'd85, 8'd93, 8'd113, 8'd115, 8'd167, 8'd95, 8'd72, 8'd139, 8'd150, 8'd125, 8'd85, 8'd119, 8'd125, 8'd93, 8'd94, 8'd169, 8'd140, 8'd154, 8'd126, 8'd150, 8'd162, 8'd118, 8'd122, 8'd184, 8'd117, 8'd116, 8'd154, 8'd94, 8'd117, 8'd184, 8'd113, 8'd100, 8'd73, 8'd142, 8'd157, 8'd111, 8'd135, 8'd52, 8'd89, 8'd129, 8'd57, 8'd125, 8'd68, 8'd132, 8'd146, 8'd145, 8'd151, 8'd170, 8'd137, 8'd119, 8'd157, 8'd154, 8'd103, 8'd184, 8'd127, 8'd114, 8'd169, 8'd198, 8'd106, 8'd71, 8'd135, 8'd109, 8'd123, 8'd84, 8'd109, 8'd58, 8'd50, 8'd82, 8'd91, 8'd66, 8'd79, 8'd95, 8'd138, 8'd164, 8'd140, 8'd189, 8'd184, 8'd134, 8'd119, 8'd134, 8'd95, 8'd171, 8'd113, 8'd154, 8'd160, 8'd179, 8'd94, 8'd102, 8'd155, 8'd78, 8'd107, 8'd82, 8'd57, 8'd98, 8'd87, 8'd103, 8'd76, 8'd150, 8'd96, 8'd160, 8'd122, 8'd150, 8'd105, 8'd85, 8'd91, 8'd87, 8'd141, 8'd151, 8'd164, 8'd137, 8'd82, 8'd73, 8'd117, 8'd108, 8'd159, 8'd84, 8'd141, 8'd139, 8'd144, 8'd95, 8'd75, 8'd78, 8'd65, 8'd101, 8'd78, 8'd120, 8'd106, 8'd99, 8'd127, 8'd162, 8'd86, 8'd150, 8'd94, 8'd140, 8'd153, 8'd139, 8'd112, 8'd133, 8'd154, 8'd138, 8'd106, 8'd113, 8'd80, 8'd99, 8'd148, 8'd110, 8'd125, 8'd101, 8'd107, 8'd132, 8'd149, 8'd123, 8'd61, 8'd107, 8'd102, 8'd147, 8'd156, 8'd79, 8'd164, 8'd103, 8'd161, 8'd128, 8'd147, 8'd138, 8'd165, 8'd94, 8'd101, 8'd155, 8'd134, 8'd180, 8'd140, 8'd172, 8'd86, 8'd120, 8'd109, 8'd95, 8'd127, 8'd140, 8'd94, 8'd149, 8'd115, 8'd145, 8'd146, 8'd143, 8'd129, 8'd93, 8'd127, 8'd75, 8'd131, 8'd150, 8'd110, 8'd141, 8'd133, 8'd114, 8'd130, 8'd93, 8'd97, 8'd161, 8'd182, 8'd134, 8'd90, 8'd106, 8'd108, 8'd44, 8'd117, 8'd142, 8'd150, 8'd126, 8'd120, 8'd81, 8'd137, 8'd106, 8'd122, 8'd83, 8'd101, 8'd97, 8'd118, 8'd119, 8'd49, 8'd75, 8'd90, 8'd124, 8'd107, 8'd94, 8'd174, 8'd182, 8'd168, 8'd152, 8'd122, 8'd86, 8'd137, 8'd111, 8'd100, 8'd109, 8'd86, 8'd111, 8'd102, 8'd154, 8'd163, 8'd121, 8'd96, 8'd90, 8'd87, 8'd99, 8'd30, 8'd106, 8'd97, 8'd84, 8'd133, 8'd105, 8'd136, 8'd88, 8'd132, 8'd116, 8'd89, 8'd134, 8'd148, 8'd92, 8'd48, 8'd90, 8'd132, 8'd116, 8'd118, 8'd109, 8'd111, 8'd126, 8'd145, 8'd81, 8'd77, 8'd52, 8'd105, 8'd95, 8'd55, 8'd130, 8'd117, 8'd101, 8'd67, 8'd156, 8'd79, 8'd128, 8'd104, 8'd102, 8'd157, 8'd115, 8'd98, 8'd145, 8'd52, 8'd106, 8'd162, 8'd129, 8'd166, 8'd152, 8'd168, 8'd133, 8'd170, 8'd101, 8'd143, 8'd60, 8'd114, 8'd72, 8'd101, 8'd106, 8'd156, 8'd79, 8'd78, 8'd147, 8'd71, 8'd150, 8'd111, 8'd147, 8'd143, 8'd170, 8'd89, 8'd83, 8'd45, 8'd85, 8'd175, 8'd154, 8'd125, 8'd160, 8'd101, 8'd169, 8'd163, 8'd138, 8'd59, 8'd60, 8'd86, 8'd105, 8'd136, 8'd57, 8'd64, 8'd150, 8'd78, 8'd129, 8'd163, 8'd162, 8'd108, 8'd125, 8'd157, 8'd91, 8'd96, 8'd88, 8'd100, 8'd103, 8'd158, 8'd141, 8'd114, 8'd153, 8'd140, 8'd157, 8'd165, 8'd82, 8'd76, 8'd69, 8'd62, 8'd146, 8'd117, 8'd104, 8'd161, 8'd127, 8'd127, 8'd162, 8'd123, 8'd188, 8'd166, 8'd134, 8'd139, 8'd163, 8'd164, 8'd170, 8'd141, 8'd122, 8'd129, 8'd146, 8'd84, 8'd143, 8'd124, 8'd97, 8'd96, 8'd145, 8'd138, 8'd79, 8'd90, 8'd166, 8'd106, 8'd127, 8'd84, 8'd143, 8'd122, 8'd167, 8'd102, 8'd165, 8'd171, 8'd161, 8'd193, 8'd169, 8'd139, 8'd150, 8'd133, 8'd146, 8'd128, 8'd132, 8'd109, 8'd134, 8'd94, 8'd90, 8'd183, 8'd145, 8'd161, 8'd107, 8'd127, 8'd141, 8'd109, 8'd109, 8'd120, 8'd78, 8'd97, 8'd156, 8'd124, 8'd142, 8'd141, 8'd130, 8'd114, 8'd186, 8'd143, 8'd127, 8'd144, 8'd199, 8'd209, 8'd160, 8'd170, 8'd122, 8'd110, 8'd161, 8'd173, 8'd153, 8'd115, 8'd135, 8'd126, 8'd190, 8'd147, 8'd155, 8'd98, 8'd143, 8'd70, 8'd111, 8'd118, 8'd110, 8'd148, 8'd174, 8'd101, 8'd88, 8'd97, 8'd96, 8'd124, 8'd161, 8'd202, 8'd138, 8'd133, 8'd126, 8'd167, 8'd112, 8'd162, 8'd179, 8'd131, 8'd159, 8'd106, 8'd117, 8'd139, 8'd131, 8'd85, 8'd158, 8'd133, 8'd98, 8'd136, 8'd78, 8'd140, 8'd181, 8'd175, 8'd169, 8'd168, 8'd94, 8'd117, 8'd174, 8'd115, 8'd136, 8'd95, 8'd132, 8'd179, 8'd102, 8'd102, 8'd155, 8'd99, 8'd100, 8'd176, 8'd112, 8'd94, 8'd109, 8'd167, 8'd111, 8'd75, 8'd168, 8'd126, 8'd123, 8'd88, 8'd109, 8'd100, 8'd109, 8'd158, 8'd135, 8'd83, 8'd82, 8'd98, 8'd136, 8'd158, 8'd116, 8'd113, 8'd130, 8'd172, 8'd182, 8'd156, 8'd131, 8'd113, 8'd116, 8'd110, 8'd174, 8'd101, 8'd145, 8'd169, 8'd163, 8'd155, 8'd104, 8'd156, 8'd104, 8'd86, 8'd118, 8'd144, 8'd117, 8'd105, 8'd100, 8'd116, 8'd72, 8'd151, 8'd95, 8'd116, 8'd146, 8'd158, 8'd107, 8'd144, 8'd159, 8'd103, 8'd107, 8'd84, 8'd143, 8'd81, 8'd136, 8'd122, 8'd82, 8'd175, 8'd158, 8'd109, 8'd139, 8'd149, 8'd161, 8'd106, 8'd125, 8'd112, 8'd141, 8'd107, 8'd93, 8'd80, 8'd121, 8'd72, 8'd146, 8'd69, 8'd124, 8'd105, 8'd117, 8'd150, 8'd117, 8'd154, 8'd135, 8'd120, 8'd112, 8'd138, 8'd110, 8'd96, 8'd71, 8'd103, 8'd87, 8'd72, 8'd144, 8'd85, 8'd77, 8'd145, 8'd107, 8'd160, 8'd136, 8'd87, 8'd112, 8'd103, 8'd84, 8'd143, 8'd151, 8'd157, 8'd154, 8'd119, 8'd103, 8'd89, 8'd152, 8'd134, 8'd129, 8'd99, 8'd136, 8'd161, 8'd137, 8'd170, 8'd110, 8'd101, 8'd121, 8'd104, 8'd109, 8'd170, 8'd107, 8'd89, 8'd131, 8'd173, 8'd141, 8'd167, 8'd164, 8'd177, 8'd167, 8'd82, 8'd152, 8'd167, 8'd130, 8'd72, 8'd113, 8'd118, 8'd145, 8'd151, 8'd106, 8'd95, 8'd84, 8'd154, 8'd115, 8'd120, 8'd95, 8'd164, 8'd120, 8'd158, 8'd163, 8'd75, 8'd102, 8'd160, 8'd140, 8'd103, 8'd111, 8'd105, 8'd148, 8'd139, 8'd108, 8'd79, 8'd123, 8'd133, 8'd175, 8'd175, 8'd104, 8'd150, 8'd112, 8'd98, 8'd127, 8'd131, 8'd92, 8'd73, 8'd78, 8'd130, 8'd103, 8'd131, 8'd73, 8'd90, 8'd109, 8'd154, 8'd137, 8'd125, 8'd109, 8'd98, 8'd87, 8'd114, 8'd137, 8'd103, 8'd164, 8'd130, 8'd132, 8'd179, 8'd185, 8'd117, 8'd125, 8'd183, 8'd142, 8'd167, 8'd70, 8'd95, 8'd100, 8'd79, 8'd93, 8'd127, 8'd155, 8'd112, 8'd145, 8'd128, 8'd162, 8'd101, 8'd125, 8'd145, 8'd112, 8'd99, 8'd159, 8'd100, 8'd108, 8'd119, 8'd145, 8'd85, 8'd109, 8'd74, 8'd73, 8'd131, 8'd157, 8'd103, 8'd149, 8'd75, 8'd131, 8'd114})
) cell_0_99 (
    .clk(clk),
    .input_index(index_0_98_99),
    .input_value(value_0_98_99),
    .input_result(result_0_98_99),
    .input_enable(enable_0_98_99),
    .output_index(index_0_99_100),
    .output_value(value_0_99_100),
    .output_result(result_0_99_100),
    .output_enable(enable_0_99_100)
);

wire [7-1:0] scale_index_0;
wire [`DATA_WIDTH-1:0] scale_value_0;
wire scale_enable_0;
scaler #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(7),
    .SCALING_FACTOR(1265583718),
    .SHIFT_AMOUNT(43),
    .OUTPUT_OFFSET(121),
    .CELL_AMOUNT(100)
) scaler_0 (
    .clk(clk),
    .input_result(result_0_99_100),
    .output_index(scale_index_0),
    .output_value(scale_value_0),
    .output_enable(scale_enable_0)
);

wire [7-1:0] index_1_0_1;
wire [`DATA_WIDTH-1:0] value_1_0_1;
wire [`DATA_WIDTH*4:0] result_1_0_1;
wire enable_1_0_1;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(7),
    .WEIGHT_AMOUNT(100),
    .WEIGHT_OFFSET(123),
    .INPUT_OFFSET(121),
    .WEIGHTS({8'd96, 8'd34, 8'd103, 8'd158, 8'd211, 8'd89, 8'd57, 8'd212, 8'd115, 8'd207, 8'd174, 8'd205, 8'd71, 8'd45, 8'd68, 8'd192, 8'd90, 8'd50, 8'd194, 8'd82, 8'd98, 8'd97, 8'd202, 8'd78, 8'd218, 8'd107, 8'd223, 8'd146, 8'd207, 8'd95, 8'd202, 8'd99, 8'd82, 8'd61, 8'd192, 8'd54, 8'd60, 8'd92, 8'd101, 8'd181, 8'd159, 8'd43, 8'd44, 8'd150, 8'd126, 8'd18, 8'd185, 8'd33, 8'd66, 8'd180, 8'd210, 8'd147, 8'd88, 8'd43, 8'd119, 8'd57, 8'd86, 8'd77, 8'd54, 8'd68, 8'd171, 8'd123, 8'd61, 8'd110, 8'd154, 8'd102, 8'd179, 8'd189, 8'd197, 8'd151, 8'd165, 8'd74, 8'd74, 8'd208, 8'd191, 8'd89, 8'd192, 8'd221, 8'd38, 8'd134, 8'd135, 8'd154, 8'd140, 8'd70, 8'd115, 8'd67, 8'd71, 8'd62, 8'd162, 8'd65, 8'd183, 8'd198, 8'd180, 8'd96, 8'd124, 8'd205, 8'd100, 8'd92, 8'd69, 8'd143})
) cell_1_0 (
    .clk(clk),
    .input_index(scale_index_0),
    .input_value(scale_value_0),
    .input_result(ground),
    .input_enable(scale_enable_0),
    .output_index(index_1_0_1),
    .output_value(value_1_0_1),
    .output_result(result_1_0_1),
    .output_enable(enable_1_0_1)
);

wire [7-1:0] index_1_1_2;
wire [`DATA_WIDTH-1:0] value_1_1_2;
wire [`DATA_WIDTH*4:0] result_1_1_2;
wire enable_1_1_2;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(7),
    .WEIGHT_AMOUNT(100),
    .WEIGHT_OFFSET(123),
    .INPUT_OFFSET(121),
    .WEIGHTS({8'd152, 8'd107, 8'd92, 8'd60, 8'd58, 8'd222, 8'd216, 8'd109, 8'd130, 8'd66, 8'd199, 8'd111, 8'd109, 8'd132, 8'd131, 8'd109, 8'd134, 8'd59, 8'd123, 8'd38, 8'd187, 8'd207, 8'd189, 8'd200, 8'd78, 8'd160, 8'd115, 8'd52, 8'd75, 8'd163, 8'd65, 8'd3, 8'd134, 8'd203, 8'd110, 8'd176, 8'd176, 8'd183, 8'd97, 8'd21, 8'd152, 8'd23, 8'd126, 8'd57, 8'd222, 8'd43, 8'd224, 8'd174, 8'd221, 8'd242, 8'd176, 8'd22, 8'd109, 8'd147, 8'd178, 8'd171, 8'd131, 8'd160, 8'd143, 8'd76, 8'd219, 8'd238, 8'd186, 8'd140, 8'd215, 8'd185, 8'd200, 8'd139, 8'd67, 8'd214, 8'd31, 8'd224, 8'd165, 8'd72, 8'd87, 8'd71, 8'd203, 8'd197, 8'd49, 8'd80, 8'd41, 8'd71, 8'd55, 8'd179, 8'd225, 8'd174, 8'd163, 8'd158, 8'd178, 8'd98, 8'd99, 8'd141, 8'd151, 8'd173, 8'd137, 8'd147, 8'd14, 8'd137, 8'd151, 8'd79})
) cell_1_1 (
    .clk(clk),
    .input_index(index_1_0_1),
    .input_value(value_1_0_1),
    .input_result(result_1_0_1),
    .input_enable(enable_1_0_1),
    .output_index(index_1_1_2),
    .output_value(value_1_1_2),
    .output_result(result_1_1_2),
    .output_enable(enable_1_1_2)
);

wire [7-1:0] index_1_2_3;
wire [`DATA_WIDTH-1:0] value_1_2_3;
wire [`DATA_WIDTH*4:0] result_1_2_3;
wire enable_1_2_3;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(7),
    .WEIGHT_AMOUNT(100),
    .WEIGHT_OFFSET(123),
    .INPUT_OFFSET(121),
    .WEIGHTS({8'd77, 8'd176, 8'd138, 8'd48, 8'd200, 8'd80, 8'd101, 8'd143, 8'd170, 8'd204, 8'd90, 8'd145, 8'd26, 8'd169, 8'd80, 8'd105, 8'd159, 8'd63, 8'd48, 8'd104, 8'd41, 8'd134, 8'd44, 8'd46, 8'd255, 8'd194, 8'd220, 8'd122, 8'd206, 8'd89, 8'd170, 8'd213, 8'd44, 8'd70, 8'd32, 8'd57, 8'd190, 8'd38, 8'd111, 8'd110, 8'd18, 8'd45, 8'd202, 8'd93, 8'd154, 8'd61, 8'd56, 8'd216, 8'd51, 8'd149, 8'd91, 8'd91, 8'd198, 8'd84, 8'd95, 8'd155, 8'd204, 8'd105, 8'd163, 8'd143, 8'd18, 8'd41, 8'd184, 8'd168, 8'd218, 8'd226, 8'd188, 8'd68, 8'd119, 8'd61, 8'd138, 8'd105, 8'd195, 8'd171, 8'd244, 8'd180, 8'd78, 8'd185, 8'd43, 8'd46, 8'd135, 8'd170, 8'd133, 8'd219, 8'd209, 8'd163, 8'd179, 8'd141, 8'd152, 8'd208, 8'd59, 8'd78, 8'd92, 8'd147, 8'd204, 8'd72, 8'd158, 8'd195, 8'd101, 8'd79})
) cell_1_2 (
    .clk(clk),
    .input_index(index_1_1_2),
    .input_value(value_1_1_2),
    .input_result(result_1_1_2),
    .input_enable(enable_1_1_2),
    .output_index(index_1_2_3),
    .output_value(value_1_2_3),
    .output_result(result_1_2_3),
    .output_enable(enable_1_2_3)
);

wire [7-1:0] index_1_3_4;
wire [`DATA_WIDTH-1:0] value_1_3_4;
wire [`DATA_WIDTH*4:0] result_1_3_4;
wire enable_1_3_4;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(7),
    .WEIGHT_AMOUNT(100),
    .WEIGHT_OFFSET(123),
    .INPUT_OFFSET(121),
    .WEIGHTS({8'd93, 8'd90, 8'd214, 8'd199, 8'd224, 8'd169, 8'd80, 8'd182, 8'd83, 8'd90, 8'd58, 8'd198, 8'd201, 8'd108, 8'd41, 8'd227, 8'd224, 8'd107, 8'd162, 8'd190, 8'd140, 8'd161, 8'd95, 8'd38, 8'd204, 8'd58, 8'd149, 8'd44, 8'd43, 8'd123, 8'd109, 8'd62, 8'd102, 8'd208, 8'd121, 8'd155, 8'd97, 8'd152, 8'd132, 8'd209, 8'd145, 8'd145, 8'd165, 8'd199, 8'd134, 8'd29, 8'd91, 8'd31, 8'd214, 8'd98, 8'd174, 8'd109, 8'd86, 8'd213, 8'd105, 8'd155, 8'd32, 8'd185, 8'd21, 8'd101, 8'd121, 8'd192, 8'd166, 8'd174, 8'd95, 8'd66, 8'd137, 8'd133, 8'd112, 8'd120, 8'd105, 8'd89, 8'd153, 8'd80, 8'd208, 8'd141, 8'd138, 8'd68, 8'd91, 8'd166, 8'd39, 8'd65, 8'd46, 8'd36, 8'd98, 8'd198, 8'd54, 8'd168, 8'd23, 8'd59, 8'd172, 8'd158, 8'd213, 8'd89, 8'd158, 8'd161, 8'd61, 8'd224, 8'd153, 8'd204})
) cell_1_3 (
    .clk(clk),
    .input_index(index_1_2_3),
    .input_value(value_1_2_3),
    .input_result(result_1_2_3),
    .input_enable(enable_1_2_3),
    .output_index(index_1_3_4),
    .output_value(value_1_3_4),
    .output_result(result_1_3_4),
    .output_enable(enable_1_3_4)
);

wire [7-1:0] index_1_4_5;
wire [`DATA_WIDTH-1:0] value_1_4_5;
wire [`DATA_WIDTH*4:0] result_1_4_5;
wire enable_1_4_5;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(7),
    .WEIGHT_AMOUNT(100),
    .WEIGHT_OFFSET(123),
    .INPUT_OFFSET(121),
    .WEIGHTS({8'd123, 8'd57, 8'd52, 8'd47, 8'd69, 8'd188, 8'd170, 8'd174, 8'd87, 8'd177, 8'd67, 8'd116, 8'd89, 8'd142, 8'd171, 8'd143, 8'd158, 8'd184, 8'd126, 8'd68, 8'd199, 8'd119, 8'd197, 8'd81, 8'd66, 8'd34, 8'd153, 8'd205, 8'd70, 8'd109, 8'd99, 8'd123, 8'd183, 8'd48, 8'd44, 8'd34, 8'd212, 8'd88, 8'd74, 8'd165, 8'd117, 8'd205, 8'd202, 8'd183, 8'd44, 8'd134, 8'd46, 8'd96, 8'd184, 8'd189, 8'd164, 8'd181, 8'd168, 8'd144, 8'd135, 8'd177, 8'd92, 8'd128, 8'd196, 8'd214, 8'd157, 8'd199, 8'd71, 8'd141, 8'd197, 8'd110, 8'd138, 8'd218, 8'd183, 8'd33, 8'd53, 8'd105, 8'd160, 8'd143, 8'd176, 8'd32, 8'd181, 8'd64, 8'd60, 8'd57, 8'd137, 8'd100, 8'd115, 8'd106, 8'd181, 8'd57, 8'd50, 8'd165, 8'd135, 8'd131, 8'd103, 8'd67, 8'd84, 8'd203, 8'd202, 8'd31, 8'd31, 8'd147, 8'd223, 8'd43})
) cell_1_4 (
    .clk(clk),
    .input_index(index_1_3_4),
    .input_value(value_1_3_4),
    .input_result(result_1_3_4),
    .input_enable(enable_1_3_4),
    .output_index(index_1_4_5),
    .output_value(value_1_4_5),
    .output_result(result_1_4_5),
    .output_enable(enable_1_4_5)
);

wire [7-1:0] index_1_5_6;
wire [`DATA_WIDTH-1:0] value_1_5_6;
wire [`DATA_WIDTH*4:0] result_1_5_6;
wire enable_1_5_6;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(7),
    .WEIGHT_AMOUNT(100),
    .WEIGHT_OFFSET(123),
    .INPUT_OFFSET(121),
    .WEIGHTS({8'd18, 8'd45, 8'd179, 8'd174, 8'd121, 8'd147, 8'd183, 8'd213, 8'd81, 8'd114, 8'd135, 8'd218, 8'd20, 8'd87, 8'd211, 8'd131, 8'd19, 8'd53, 8'd50, 8'd138, 8'd192, 8'd165, 8'd143, 8'd126, 8'd141, 8'd151, 8'd112, 8'd191, 8'd109, 8'd221, 8'd63, 8'd209, 8'd20, 8'd154, 8'd199, 8'd207, 8'd169, 8'd81, 8'd195, 8'd136, 8'd170, 8'd145, 8'd165, 8'd226, 8'd156, 8'd179, 8'd159, 8'd187, 8'd85, 8'd123, 8'd185, 8'd172, 8'd32, 8'd209, 8'd54, 8'd82, 8'd177, 8'd16, 8'd35, 8'd80, 8'd30, 8'd188, 8'd114, 8'd34, 8'd170, 8'd169, 8'd177, 8'd166, 8'd137, 8'd29, 8'd125, 8'd84, 8'd138, 8'd61, 8'd129, 8'd192, 8'd168, 8'd61, 8'd175, 8'd79, 8'd64, 8'd165, 8'd224, 8'd182, 8'd82, 8'd55, 8'd145, 8'd205, 8'd173, 8'd174, 8'd112, 8'd70, 8'd156, 8'd171, 8'd120, 8'd178, 8'd95, 8'd138, 8'd112, 8'd217})
) cell_1_5 (
    .clk(clk),
    .input_index(index_1_4_5),
    .input_value(value_1_4_5),
    .input_result(result_1_4_5),
    .input_enable(enable_1_4_5),
    .output_index(index_1_5_6),
    .output_value(value_1_5_6),
    .output_result(result_1_5_6),
    .output_enable(enable_1_5_6)
);

wire [7-1:0] index_1_6_7;
wire [`DATA_WIDTH-1:0] value_1_6_7;
wire [`DATA_WIDTH*4:0] result_1_6_7;
wire enable_1_6_7;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(7),
    .WEIGHT_AMOUNT(100),
    .WEIGHT_OFFSET(123),
    .INPUT_OFFSET(121),
    .WEIGHTS({8'd215, 8'd26, 8'd141, 8'd149, 8'd79, 8'd233, 8'd181, 8'd198, 8'd213, 8'd95, 8'd174, 8'd121, 8'd129, 8'd141, 8'd53, 8'd16, 8'd115, 8'd92, 8'd221, 8'd180, 8'd41, 8'd78, 8'd211, 8'd51, 8'd82, 8'd77, 8'd204, 8'd67, 8'd159, 8'd182, 8'd45, 8'd83, 8'd26, 8'd48, 8'd80, 8'd48, 8'd155, 8'd38, 8'd86, 8'd139, 8'd70, 8'd141, 8'd52, 8'd58, 8'd232, 8'd240, 8'd193, 8'd95, 8'd74, 8'd206, 8'd50, 8'd70, 8'd72, 8'd134, 8'd98, 8'd48, 8'd77, 8'd205, 8'd174, 8'd196, 8'd46, 8'd214, 8'd40, 8'd162, 8'd187, 8'd153, 8'd87, 8'd222, 8'd152, 8'd165, 8'd109, 8'd235, 8'd165, 8'd89, 8'd157, 8'd91, 8'd123, 8'd196, 8'd107, 8'd33, 8'd123, 8'd205, 8'd152, 8'd182, 8'd164, 8'd107, 8'd159, 8'd94, 8'd135, 8'd98, 8'd67, 8'd167, 8'd129, 8'd192, 8'd148, 8'd233, 8'd97, 8'd45, 8'd70, 8'd139})
) cell_1_6 (
    .clk(clk),
    .input_index(index_1_5_6),
    .input_value(value_1_5_6),
    .input_result(result_1_5_6),
    .input_enable(enable_1_5_6),
    .output_index(index_1_6_7),
    .output_value(value_1_6_7),
    .output_result(result_1_6_7),
    .output_enable(enable_1_6_7)
);

wire [7-1:0] index_1_7_8;
wire [`DATA_WIDTH-1:0] value_1_7_8;
wire [`DATA_WIDTH*4:0] result_1_7_8;
wire enable_1_7_8;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(7),
    .WEIGHT_AMOUNT(100),
    .WEIGHT_OFFSET(123),
    .INPUT_OFFSET(121),
    .WEIGHTS({8'd118, 8'd61, 8'd61, 8'd71, 8'd171, 8'd124, 8'd127, 8'd156, 8'd85, 8'd112, 8'd112, 8'd64, 8'd80, 8'd45, 8'd176, 8'd43, 8'd48, 8'd56, 8'd195, 8'd167, 8'd205, 8'd81, 8'd135, 8'd114, 8'd46, 8'd74, 8'd184, 8'd201, 8'd73, 8'd208, 8'd206, 8'd45, 8'd100, 8'd86, 8'd95, 8'd92, 8'd94, 8'd207, 8'd109, 8'd103, 8'd102, 8'd113, 8'd69, 8'd77, 8'd128, 8'd139, 8'd200, 8'd154, 8'd164, 8'd150, 8'd65, 8'd111, 8'd88, 8'd84, 8'd189, 8'd38, 8'd202, 8'd182, 8'd104, 8'd78, 8'd108, 8'd109, 8'd157, 8'd94, 8'd219, 8'd37, 8'd61, 8'd205, 8'd124, 8'd180, 8'd162, 8'd44, 8'd144, 8'd155, 8'd45, 8'd23, 8'd149, 8'd65, 8'd151, 8'd194, 8'd117, 8'd95, 8'd186, 8'd82, 8'd150, 8'd35, 8'd114, 8'd136, 8'd56, 8'd77, 8'd158, 8'd137, 8'd153, 8'd61, 8'd54, 8'd61, 8'd86, 8'd89, 8'd192, 8'd137})
) cell_1_7 (
    .clk(clk),
    .input_index(index_1_6_7),
    .input_value(value_1_6_7),
    .input_result(result_1_6_7),
    .input_enable(enable_1_6_7),
    .output_index(index_1_7_8),
    .output_value(value_1_7_8),
    .output_result(result_1_7_8),
    .output_enable(enable_1_7_8)
);

wire [7-1:0] index_1_8_9;
wire [`DATA_WIDTH-1:0] value_1_8_9;
wire [`DATA_WIDTH*4:0] result_1_8_9;
wire enable_1_8_9;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(7),
    .WEIGHT_AMOUNT(100),
    .WEIGHT_OFFSET(123),
    .INPUT_OFFSET(121),
    .WEIGHTS({8'd76, 8'd29, 8'd37, 8'd12, 8'd4, 8'd151, 8'd53, 8'd144, 8'd190, 8'd111, 8'd10, 8'd132, 8'd125, 8'd169, 8'd128, 8'd201, 8'd101, 8'd91, 8'd81, 8'd202, 8'd222, 8'd171, 8'd173, 8'd24, 8'd48, 8'd70, 8'd180, 8'd195, 8'd162, 8'd113, 8'd30, 8'd166, 8'd145, 8'd68, 8'd83, 8'd211, 8'd59, 8'd83, 8'd83, 8'd110, 8'd41, 8'd60, 8'd99, 8'd53, 8'd216, 8'd129, 8'd188, 8'd124, 8'd142, 8'd199, 8'd39, 8'd33, 8'd200, 8'd144, 8'd110, 8'd134, 8'd202, 8'd61, 8'd85, 8'd24, 8'd108, 8'd211, 8'd96, 8'd109, 8'd170, 8'd31, 8'd120, 8'd29, 8'd56, 8'd215, 8'd81, 8'd174, 8'd215, 8'd202, 8'd49, 8'd221, 8'd82, 8'd199, 8'd156, 8'd53, 8'd129, 8'd94, 8'd67, 8'd84, 8'd117, 8'd30, 8'd57, 8'd208, 8'd14, 8'd79, 8'd204, 8'd215, 8'd152, 8'd156, 8'd128, 8'd97, 8'd83, 8'd225, 8'd53, 8'd124})
) cell_1_8 (
    .clk(clk),
    .input_index(index_1_7_8),
    .input_value(value_1_7_8),
    .input_result(result_1_7_8),
    .input_enable(enable_1_7_8),
    .output_index(index_1_8_9),
    .output_value(value_1_8_9),
    .output_result(result_1_8_9),
    .output_enable(enable_1_8_9)
);

wire [7-1:0] index_1_9_10;
wire [`DATA_WIDTH-1:0] value_1_9_10;
wire [`DATA_WIDTH*4:0] result_1_9_10;
wire enable_1_9_10;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(7),
    .WEIGHT_AMOUNT(100),
    .WEIGHT_OFFSET(123),
    .INPUT_OFFSET(121),
    .WEIGHTS({8'd148, 8'd161, 8'd90, 8'd160, 8'd164, 8'd192, 8'd124, 8'd68, 8'd89, 8'd42, 8'd103, 8'd42, 8'd29, 8'd203, 8'd114, 8'd134, 8'd46, 8'd183, 8'd92, 8'd162, 8'd103, 8'd144, 8'd204, 8'd149, 8'd171, 8'd177, 8'd175, 8'd138, 8'd90, 8'd153, 8'd185, 8'd149, 8'd130, 8'd179, 8'd37, 8'd137, 8'd85, 8'd63, 8'd27, 8'd61, 8'd37, 8'd31, 8'd224, 8'd198, 8'd60, 8'd30, 8'd161, 8'd89, 8'd157, 8'd37, 8'd109, 8'd81, 8'd82, 8'd149, 8'd148, 8'd194, 8'd152, 8'd97, 8'd41, 8'd141, 8'd66, 8'd87, 8'd78, 8'd176, 8'd158, 8'd34, 8'd227, 8'd167, 8'd24, 8'd40, 8'd224, 8'd8, 8'd143, 8'd157, 8'd222, 8'd55, 8'd106, 8'd193, 8'd194, 8'd76, 8'd67, 8'd222, 8'd75, 8'd54, 8'd0, 8'd29, 8'd127, 8'd117, 8'd110, 8'd92, 8'd199, 8'd144, 8'd230, 8'd76, 8'd226, 8'd105, 8'd53, 8'd93, 8'd72, 8'd169})
) cell_1_9 (
    .clk(clk),
    .input_index(index_1_8_9),
    .input_value(value_1_8_9),
    .input_result(result_1_8_9),
    .input_enable(enable_1_8_9),
    .output_index(index_1_9_10),
    .output_value(value_1_9_10),
    .output_result(result_1_9_10),
    .output_enable(enable_1_9_10)
);

wire [4-1:0] scale_index_1;
wire [`DATA_WIDTH-1:0] scale_value_1;
wire scale_enable_1;
scaler #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(4),
    .SCALING_FACTOR(1960168069),
    .SHIFT_AMOUNT(41),
    .OUTPUT_OFFSET(127),
    .CELL_AMOUNT(10)
) scaler_1 (
    .clk(clk),
    .input_result(result_1_9_10),
    .output_index(scale_index_1),
    .output_value(scale_value_1),
    .output_enable(scale_enable_1)
);

wire [4-1:0] index_2_0_1;
wire [`DATA_WIDTH-1:0] value_2_0_1;
wire [`DATA_WIDTH*4:0] result_2_0_1;
wire enable_2_0_1;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(4),
    .WEIGHT_AMOUNT(10),
    .WEIGHT_OFFSET(127),
    .INPUT_OFFSET(127),
    .WEIGHTS({8'd170, 8'd127, 8'd153, 8'd140, 8'd9, 8'd221, 8'd224, 8'd24, 8'd183, 8'd56})
) cell_2_0 (
    .clk(clk),
    .input_index(scale_index_1),
    .input_value(scale_value_1),
    .input_result(ground),
    .input_enable(scale_enable_1),
    .output_index(index_2_0_1),
    .output_value(value_2_0_1),
    .output_result(result_2_0_1),
    .output_enable(enable_2_0_1)
);

wire [4-1:0] index_2_1_2;
wire [`DATA_WIDTH-1:0] value_2_1_2;
wire [`DATA_WIDTH*4:0] result_2_1_2;
wire enable_2_1_2;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(4),
    .WEIGHT_AMOUNT(10),
    .WEIGHT_OFFSET(127),
    .INPUT_OFFSET(127),
    .WEIGHTS({8'd130, 8'd171, 8'd21, 8'd231, 8'd196, 8'd212, 8'd113, 8'd198, 8'd93, 8'd77})
) cell_2_1 (
    .clk(clk),
    .input_index(index_2_0_1),
    .input_value(value_2_0_1),
    .input_result(result_2_0_1),
    .input_enable(enable_2_0_1),
    .output_index(index_2_1_2),
    .output_value(value_2_1_2),
    .output_result(result_2_1_2),
    .output_enable(enable_2_1_2)
);

wire [4-1:0] index_2_2_3;
wire [`DATA_WIDTH-1:0] value_2_2_3;
wire [`DATA_WIDTH*4:0] result_2_2_3;
wire enable_2_2_3;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(4),
    .WEIGHT_AMOUNT(10),
    .WEIGHT_OFFSET(127),
    .INPUT_OFFSET(127),
    .WEIGHTS({8'd150, 8'd228, 8'd231, 8'd53, 8'd213, 8'd157, 8'd100, 8'd93, 8'd216, 8'd118})
) cell_2_2 (
    .clk(clk),
    .input_index(index_2_1_2),
    .input_value(value_2_1_2),
    .input_result(result_2_1_2),
    .input_enable(enable_2_1_2),
    .output_index(index_2_2_3),
    .output_value(value_2_2_3),
    .output_result(result_2_2_3),
    .output_enable(enable_2_2_3)
);

wire [4-1:0] index_2_3_4;
wire [`DATA_WIDTH-1:0] value_2_3_4;
wire [`DATA_WIDTH*4:0] result_2_3_4;
wire enable_2_3_4;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(4),
    .WEIGHT_AMOUNT(10),
    .WEIGHT_OFFSET(127),
    .INPUT_OFFSET(127),
    .WEIGHTS({8'd195, 8'd158, 8'd117, 8'd250, 8'd190, 8'd128, 8'd83, 8'd16, 8'd154, 8'd105})
) cell_2_3 (
    .clk(clk),
    .input_index(index_2_2_3),
    .input_value(value_2_2_3),
    .input_result(result_2_2_3),
    .input_enable(enable_2_2_3),
    .output_index(index_2_3_4),
    .output_value(value_2_3_4),
    .output_result(result_2_3_4),
    .output_enable(enable_2_3_4)
);

wire [4-1:0] index_2_4_5;
wire [`DATA_WIDTH-1:0] value_2_4_5;
wire [`DATA_WIDTH*4:0] result_2_4_5;
wire enable_2_4_5;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(4),
    .WEIGHT_AMOUNT(10),
    .WEIGHT_OFFSET(127),
    .INPUT_OFFSET(127),
    .WEIGHTS({8'd142, 8'd118, 8'd184, 8'd41, 8'd226, 8'd81, 8'd49, 8'd33, 8'd23, 8'd134})
) cell_2_4 (
    .clk(clk),
    .input_index(index_2_3_4),
    .input_value(value_2_3_4),
    .input_result(result_2_3_4),
    .input_enable(enable_2_3_4),
    .output_index(index_2_4_5),
    .output_value(value_2_4_5),
    .output_result(result_2_4_5),
    .output_enable(enable_2_4_5)
);

wire [4-1:0] index_2_5_6;
wire [`DATA_WIDTH-1:0] value_2_5_6;
wire [`DATA_WIDTH*4:0] result_2_5_6;
wire enable_2_5_6;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(4),
    .WEIGHT_AMOUNT(10),
    .WEIGHT_OFFSET(127),
    .INPUT_OFFSET(127),
    .WEIGHTS({8'd190, 8'd45, 8'd170, 8'd165, 8'd102, 8'd50, 8'd174, 8'd55, 8'd220, 8'd255})
) cell_2_5 (
    .clk(clk),
    .input_index(index_2_4_5),
    .input_value(value_2_4_5),
    .input_result(result_2_4_5),
    .input_enable(enable_2_4_5),
    .output_index(index_2_5_6),
    .output_value(value_2_5_6),
    .output_result(result_2_5_6),
    .output_enable(enable_2_5_6)
);

wire [4-1:0] index_2_6_7;
wire [`DATA_WIDTH-1:0] value_2_6_7;
wire [`DATA_WIDTH*4:0] result_2_6_7;
wire enable_2_6_7;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(4),
    .WEIGHT_AMOUNT(10),
    .WEIGHT_OFFSET(127),
    .INPUT_OFFSET(127),
    .WEIGHTS({8'd177, 8'd185, 8'd28, 8'd100, 8'd124, 8'd95, 8'd189, 8'd64, 8'd134, 8'd39})
) cell_2_6 (
    .clk(clk),
    .input_index(index_2_5_6),
    .input_value(value_2_5_6),
    .input_result(result_2_5_6),
    .input_enable(enable_2_5_6),
    .output_index(index_2_6_7),
    .output_value(value_2_6_7),
    .output_result(result_2_6_7),
    .output_enable(enable_2_6_7)
);

wire [4-1:0] index_2_7_8;
wire [`DATA_WIDTH-1:0] value_2_7_8;
wire [`DATA_WIDTH*4:0] result_2_7_8;
wire enable_2_7_8;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(4),
    .WEIGHT_AMOUNT(10),
    .WEIGHT_OFFSET(127),
    .INPUT_OFFSET(127),
    .WEIGHTS({8'd94, 8'd108, 8'd97, 8'd123, 8'd43, 8'd82, 8'd21, 8'd96, 8'd171, 8'd54})
) cell_2_7 (
    .clk(clk),
    .input_index(index_2_6_7),
    .input_value(value_2_6_7),
    .input_result(result_2_6_7),
    .input_enable(enable_2_6_7),
    .output_index(index_2_7_8),
    .output_value(value_2_7_8),
    .output_result(result_2_7_8),
    .output_enable(enable_2_7_8)
);

wire [4-1:0] index_2_8_9;
wire [`DATA_WIDTH-1:0] value_2_8_9;
wire [`DATA_WIDTH*4:0] result_2_8_9;
wire enable_2_8_9;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(4),
    .WEIGHT_AMOUNT(10),
    .WEIGHT_OFFSET(127),
    .INPUT_OFFSET(127),
    .WEIGHTS({8'd186, 8'd54, 8'd132, 8'd106, 8'd174, 8'd225, 8'd185, 8'd158, 8'd220, 8'd81})
) cell_2_8 (
    .clk(clk),
    .input_index(index_2_7_8),
    .input_value(value_2_7_8),
    .input_result(result_2_7_8),
    .input_enable(enable_2_7_8),
    .output_index(index_2_8_9),
    .output_value(value_2_8_9),
    .output_result(result_2_8_9),
    .output_enable(enable_2_8_9)
);

wire [4-1:0] index_2_9_10;
wire [`DATA_WIDTH-1:0] value_2_9_10;
wire [`DATA_WIDTH*4:0] result_2_9_10;
wire enable_2_9_10;
weight_comp_cell #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(4),
    .WEIGHT_AMOUNT(10),
    .WEIGHT_OFFSET(127),
    .INPUT_OFFSET(127),
    .WEIGHTS({8'd0, 8'd31, 8'd128, 8'd58, 8'd195, 8'd203, 8'd193, 8'd90, 8'd181, 8'd62})
) cell_2_9 (
    .clk(clk),
    .input_index(index_2_8_9),
    .input_value(value_2_8_9),
    .input_result(result_2_8_9),
    .input_enable(enable_2_8_9),
    .output_index(index_2_9_10),
    .output_value(value_2_9_10),
    .output_result(result_2_9_10),
    .output_enable(enable_2_9_10)
);

wire [4-1:0] scale_index_2;
wire [`DATA_WIDTH-1:0] scale_value_2;
wire scale_enable_2;
scaler #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(4),
    .SCALING_FACTOR(1727327655),
    .SHIFT_AMOUNT(33),
    .OUTPUT_OFFSET(0),
    .CELL_AMOUNT(10)
) scaler_2 (
    .clk(clk),
    .input_result(result_2_9_10),
    .output_index(scale_index_2),
    .output_value(scale_value_2),
    .output_enable(scale_enable_2)
);

wire [`DATA_WIDTH*4:0] output_result;

argmax_cell  #(
    .DATA_WIDTH(`DATA_WIDTH),
    .RESULT_WIDTH(`DATA_WIDTH*4),
    .INDEX_WIDTH(4),
    .CELL_AMOUNT(10)
) result_cell (
    .clk(clk),
    .input_index(scale_index_2),
    .input_value(scale_value_2),
    .input_enable(scale_enable_2),
    .output_result(output_result)
);

initial begin
    clk = 1;
    forever #(`CLOCK/2) clk = !clk;
end

initial begin
    input_value = 0;
    input_index = 0;
    input_enable = 0;
    pixels_fed = 0;
    numbers_streamed = 0;
    open_data_file("/home/mbax4km4/FinalProject/MLontoFPGAs/VerilogSrc/Simulators/test_data/zero.txt");
end

reg [3:0] output_results_checked;
        
initial begin
    output_results_checked = 0;
end

//always @ (posedge clk) begin
//    if (result_0_99_100[`DATA_WIDTH*4]!=0) begin
//        #1
//        check_output(result_0_99_100[`DATA_WIDTH*4-1:0], 66019);
//        $stop;
//    end
//end 

//always @ (posedge clk) begin
//    if (scale_enable_1!=0) begin
//        #1
//        check_output(scale_value_1, 81);
//        #(`CLOCK)
//        check_output(scale_value_1, 192);
//        #(`CLOCK)
//        check_output(scale_value_1, 59);
//        #(`CLOCK)
//        check_output(scale_value_1, 144);
//        #(`CLOCK)
//        check_output(scale_value_1, 125);
//        $stop;
//    end
//end

//always @ (posedge clk) begin
//    if (scale_enable_2!=0) begin
//        #1
//        check_output(scale_value_2, 4148);
//        #(`CLOCK)
//        check_output(scale_value_2, -2306);
//        #(`CLOCK)
//        check_output(scale_value_2, 1776);
//        #(`CLOCK)
//        check_output(scale_value_2, 1334);
//        #(`CLOCK)
//        check_output(scale_value_2, -414);
//        $stop;
//    end
//end
    
always @ (posedge clk) begin #2
    if (pixels_fed!=file_lines_read) begin
        input_value <= pixel_data[pixels_fed];
        input_index <= pixels_fed;
        input_enable <= 1;
        if (pixels_fed + 1 == file_lines_read && numbers_streamed != 9) begin
            pixels_fed <= 0;
            if (numbers_streamed == 0) begin
                open_data_file("/home/mbax4km4/FinalProject/MLontoFPGAs/VerilogSrc/Simulators/test_data/one.txt");
            end
            if (numbers_streamed == 1) begin
                open_data_file("/home/mbax4km4/FinalProject/MLontoFPGAs/VerilogSrc/Simulators/test_data/two.txt");
            end
            if (numbers_streamed == 2) begin
                open_data_file("/home/mbax4km4/FinalProject/MLontoFPGAs/VerilogSrc/Simulators/test_data/three.txt");
            end
            if (numbers_streamed == 3) begin
                open_data_file("/home/mbax4km4/FinalProject/MLontoFPGAs/VerilogSrc/Simulators/test_data/four.txt");
            end
            if (numbers_streamed == 4) begin
                open_data_file("/home/mbax4km4/FinalProject/MLontoFPGAs/VerilogSrc/Simulators/test_data/five.txt");
            end
            if (numbers_streamed == 5) begin
                open_data_file("/home/mbax4km4/FinalProject/MLontoFPGAs/VerilogSrc/Simulators/test_data/six.txt");
            end                                                
            if (numbers_streamed == 6) begin
                open_data_file("/home/mbax4km4/FinalProject/MLontoFPGAs/VerilogSrc/Simulators/test_data/seven.txt");
            end
            if (numbers_streamed == 7) begin
                open_data_file("/home/mbax4km4/FinalProject/MLontoFPGAs/VerilogSrc/Simulators/test_data/eight.txt");
            end
            if (numbers_streamed == 8) begin
                open_data_file("/home/mbax4km4/FinalProject/MLontoFPGAs/VerilogSrc/Simulators/test_data/nine.txt");
            end                                         
            numbers_streamed <= numbers_streamed + 1;
        end
        else begin
            pixels_fed <= pixels_fed + 1;
        end
    end
    else begin
        input_enable <= 0;
    end
    if (output_result[`DATA_WIDTH*4]) begin
        output_results_checked <= output_results_checked+1;
        if (output_results_checked == 0) begin
            check_output(output_result[`DATA_WIDTH*4-1:0], 0);
        end
        if (output_results_checked == 1) begin
            check_output(output_result[`DATA_WIDTH*4-1:0], 1);
        end
        if (output_results_checked == 2) begin
            check_output(output_result[`DATA_WIDTH*4-1:0], 2);
        end
        if (output_results_checked == 3) begin
            check_output(output_result[`DATA_WIDTH*4-1:0], 3);
        end
        if (output_results_checked == 4) begin
            check_output(output_result[`DATA_WIDTH*4-1:0], 4);
        end
        if (output_results_checked == 5) begin
            check_output(output_result[`DATA_WIDTH*4-1:0], 5);
        end
        if (output_results_checked == 6) begin
            check_output(output_result[`DATA_WIDTH*4-1:0], 6);
        end
        if (output_results_checked == 7) begin
            check_output(output_result[`DATA_WIDTH*4-1:0], 7);
        end
        if (output_results_checked == 8) begin
            check_output(output_result[`DATA_WIDTH*4-1:0], 8);
        end                                                                
        if (output_results_checked == 9) begin
            check_output(output_result[`DATA_WIDTH*4-1:0], 9);
            #(`CLOCK*2);
            $display("SUCCESSFUL TEST!"); 
            $stop;
        end
    end
end

endmodule
